library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity tapper_sound_cpu is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of tapper_sound_cpu is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"F3",X"31",X"FF",X"83",X"ED",X"56",X"18",X"58",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"3A",X"00",X"E0",X"3A",X"41",X"80",X"3C",
		X"32",X"41",X"80",X"F1",X"FB",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"00",X"B0",X"36",X"0F",X"21",X"02",X"B0",X"36",X"F0",X"3A",X"00",X"F0",X"CB",X"47",X"20",
		X"4E",X"CB",X"4F",X"20",X"2D",X"AF",X"32",X"C7",X"81",X"CD",X"26",X"06",X"CD",X"DE",X"06",X"3A",
		X"C7",X"81",X"B7",X"28",X"1D",X"CB",X"67",X"20",X"05",X"01",X"00",X"10",X"18",X"03",X"01",X"00",
		X"80",X"11",X"01",X"00",X"60",X"69",X"32",X"00",X"D0",X"37",X"3F",X"ED",X"52",X"20",X"FC",X"2F",
		X"18",X"F2",X"3E",X"FF",X"32",X"00",X"D0",X"3A",X"00",X"F0",X"CB",X"57",X"20",X"08",X"CD",X"06",
		X"0A",X"18",X"EF",X"3A",X"00",X"F0",X"CB",X"5F",X"20",X"F9",X"CD",X"2D",X"0A",X"18",X"F4",X"06",
		X"00",X"CD",X"E9",X"09",X"06",X"FF",X"CD",X"E9",X"09",X"06",X"55",X"CD",X"E9",X"09",X"06",X"AA",
		X"CD",X"E9",X"09",X"AF",X"32",X"C7",X"81",X"CD",X"26",X"06",X"CD",X"DE",X"06",X"3A",X"C7",X"81",
		X"32",X"00",X"C0",X"CD",X"59",X"02",X"FD",X"21",X"3D",X"81",X"11",X"17",X"00",X"06",X"06",X"FD",
		X"7E",X"00",X"B7",X"28",X"4F",X"FD",X"19",X"10",X"F6",X"FD",X"21",X"3D",X"81",X"06",X"06",X"DD",
		X"7E",X"03",X"FD",X"BE",X"07",X"38",X"2D",X"FD",X"19",X"10",X"F4",X"E5",X"21",X"00",X"00",X"FD",
		X"21",X"3D",X"81",X"06",X"06",X"0E",X"10",X"FD",X"7E",X"07",X"DD",X"BE",X"03",X"20",X"0A",X"FD",
		X"7E",X"14",X"B9",X"30",X"04",X"4F",X"FD",X"E5",X"E1",X"FD",X"19",X"10",X"EA",X"7C",X"B5",X"E5",
		X"FD",X"E1",X"E1",X"C8",X"DD",X"E5",X"FD",X"56",X"06",X"FD",X"5E",X"05",X"D5",X"DD",X"E1",X"DD",
		X"35",X"18",X"DD",X"E1",X"FD",X"36",X"00",X"01",X"7E",X"FD",X"77",X"0F",X"23",X"7E",X"FD",X"77",
		X"10",X"DD",X"4E",X"06",X"23",X"5E",X"23",X"56",X"FD",X"73",X"02",X"FD",X"72",X"03",X"FD",X"71",
		X"04",X"DD",X"7E",X"03",X"FD",X"77",X"07",X"DD",X"E5",X"D1",X"FD",X"73",X"05",X"FD",X"72",X"06",
		X"AF",X"06",X"07",X"FD",X"77",X"08",X"FD",X"23",X"10",X"F9",X"DD",X"34",X"18",X"C9",X"DD",X"66",
		X"06",X"DD",X"6E",X"05",X"E5",X"FD",X"E1",X"DD",X"7E",X"00",X"DD",X"66",X"03",X"DD",X"6E",X"02",
		X"06",X"00",X"DD",X"4E",X"04",X"AF",X"ED",X"42",X"DD",X"74",X"03",X"DD",X"75",X"02",X"D0",X"FD",
		X"7E",X"01",X"FD",X"B6",X"02",X"28",X"04",X"DD",X"34",X"00",X"C9",X"DD",X"77",X"00",X"FD",X"35",
		X"18",X"CD",X"A9",X"08",X"AF",X"CD",X"C3",X"08",X"AF",X"CD",X"C3",X"08",X"C9",X"21",X"43",X"80",
		X"11",X"44",X"80",X"01",X"F9",X"00",X"36",X"00",X"ED",X"B0",X"21",X"3D",X"81",X"11",X"3E",X"81",
		X"01",X"89",X"00",X"36",X"00",X"ED",X"B0",X"DD",X"21",X"2F",X"80",X"FD",X"21",X"00",X"A0",X"21",
		X"0F",X"80",X"11",X"33",X"02",X"06",X"0F",X"1A",X"77",X"DD",X"77",X"00",X"FD",X"70",X"00",X"32",
		X"02",X"A0",X"2B",X"DD",X"2B",X"13",X"05",X"F2",X"E7",X"01",X"DD",X"21",X"3F",X"80",X"FD",X"21",
		X"00",X"B0",X"21",X"1F",X"80",X"11",X"43",X"02",X"06",X"0F",X"1A",X"77",X"DD",X"77",X"00",X"FD",
		X"70",X"00",X"32",X"02",X"B0",X"2B",X"DD",X"2B",X"13",X"05",X"F2",X"0A",X"02",X"21",X"3E",X"81",
		X"DD",X"21",X"53",X"02",X"06",X"06",X"11",X"17",X"00",X"DD",X"7E",X"00",X"77",X"19",X"DD",X"23",
		X"10",X"F7",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"01",X"04",X"02",X"05",X"31",X"FF",X"83",X"F3",X"ED",X"56",X"CD",
		X"D0",X"09",X"CD",X"D4",X"03",X"FB",X"CD",X"BF",X"03",X"CD",X"BA",X"02",X"CD",X"D4",X"03",X"21",
		X"40",X"80",X"3A",X"41",X"80",X"BE",X"38",X"FA",X"4F",X"06",X"10",X"3A",X"42",X"80",X"C6",X"40",
		X"FE",X"64",X"38",X"04",X"D6",X"64",X"06",X"0F",X"32",X"42",X"80",X"70",X"06",X"00",X"21",X"CE",
		X"81",X"09",X"34",X"AF",X"32",X"41",X"80",X"18",X"CD",X"1E",X"00",X"06",X"08",X"CB",X"7A",X"28",
		X"06",X"CB",X"3A",X"CB",X"3C",X"CB",X"1D",X"AF",X"ED",X"52",X"23",X"F2",X"B0",X"02",X"19",X"2B",
		X"29",X"10",X"F4",X"7C",X"BA",X"D8",X"2C",X"92",X"67",X"C9",X"DD",X"21",X"3D",X"81",X"06",X"06",
		X"DD",X"7E",X"00",X"B7",X"28",X"05",X"C5",X"CD",X"7E",X"01",X"C1",X"11",X"17",X"00",X"DD",X"19",
		X"10",X"EE",X"DD",X"21",X"43",X"80",X"06",X"0A",X"C5",X"DD",X"7E",X"00",X"B7",X"CA",X"60",X"03",
		X"3D",X"20",X"74",X"DD",X"66",X"05",X"DD",X"6E",X"04",X"DD",X"7E",X"06",X"CD",X"00",X"0B",X"DD",
		X"74",X"05",X"DD",X"75",X"04",X"DD",X"4E",X"16",X"DD",X"46",X"17",X"C5",X"FD",X"E1",X"FD",X"5E",
		X"00",X"FD",X"56",X"01",X"7A",X"FE",X"FF",X"20",X"33",X"DD",X"7E",X"07",X"FE",X"02",X"38",X"26",
		X"AF",X"FD",X"56",X"03",X"FD",X"5E",X"02",X"ED",X"52",X"38",X"45",X"DD",X"77",X"04",X"DD",X"77",
		X"05",X"DD",X"56",X"14",X"DD",X"5E",X"15",X"DD",X"72",X"16",X"DD",X"73",X"17",X"FE",X"FF",X"28",
		X"2F",X"DD",X"35",X"07",X"18",X"2A",X"DD",X"36",X"00",X"02",X"18",X"24",X"AF",X"ED",X"52",X"38",
		X"1F",X"FD",X"E5",X"E1",X"11",X"06",X"00",X"19",X"DD",X"74",X"17",X"DD",X"75",X"16",X"11",X"FC",
		X"FF",X"19",X"CD",X"E6",X"00",X"18",X"09",X"DD",X"7E",X"18",X"B7",X"20",X"03",X"DD",X"77",X"00",
		X"C1",X"11",X"19",X"00",X"DD",X"19",X"05",X"C2",X"D8",X"02",X"DD",X"21",X"3D",X"81",X"06",X"06",
		X"DD",X"7E",X"00",X"B7",X"28",X"05",X"C5",X"CD",X"48",X"04",X"C1",X"11",X"17",X"00",X"DD",X"19",
		X"10",X"EE",X"C9",X"DD",X"E5",X"E5",X"DD",X"E1",X"DD",X"96",X"FE",X"28",X"2C",X"67",X"0E",X"00",
		X"DD",X"7E",X"01",X"DD",X"96",X"FF",X"28",X"21",X"30",X"03",X"2F",X"3C",X"0C",X"5F",X"CD",X"09",
		X"04",X"DD",X"7E",X"00",X"DD",X"96",X"FE",X"57",X"CD",X"99",X"02",X"DD",X"7E",X"FF",X"0D",X"28",
		X"04",X"85",X"DD",X"E1",X"C9",X"95",X"DD",X"E1",X"C9",X"DD",X"7E",X"FF",X"DD",X"E1",X"C9",X"E5",
		X"21",X"C8",X"81",X"3A",X"00",X"90",X"E6",X"80",X"AE",X"28",X"07",X"7E",X"EE",X"80",X"77",X"CD",
		X"35",X"07",X"E1",X"C9",X"21",X"3F",X"80",X"11",X"1F",X"80",X"06",X"0F",X"DD",X"21",X"00",X"B0",
		X"1A",X"BE",X"28",X"07",X"77",X"DD",X"70",X"00",X"32",X"02",X"B0",X"1B",X"2B",X"05",X"F2",X"E0",
		X"03",X"06",X"0F",X"DD",X"21",X"00",X"A0",X"1A",X"BE",X"28",X"07",X"77",X"DD",X"70",X"00",X"32",
		X"02",X"A0",X"1B",X"2B",X"05",X"F2",X"F7",X"03",X"C9",X"16",X"00",X"3E",X"08",X"BC",X"30",X"0E",
		X"BB",X"30",X"0E",X"2E",X"00",X"06",X"08",X"29",X"30",X"01",X"19",X"10",X"FA",X"C9",X"44",X"18",
		X"02",X"43",X"5C",X"21",X"00",X"00",X"78",X"B7",X"C8",X"19",X"10",X"FD",X"C9",X"67",X"7A",X"B7",
		X"28",X"12",X"7C",X"06",X"10",X"21",X"00",X"00",X"CB",X"39",X"1F",X"30",X"01",X"19",X"EB",X"29",
		X"EB",X"10",X"F5",X"C9",X"CD",X"09",X"04",X"C9",X"DD",X"66",X"06",X"DD",X"6E",X"05",X"E5",X"FD",
		X"E1",X"CD",X"64",X"04",X"CD",X"F1",X"05",X"CD",X"CE",X"04",X"CD",X"5E",X"05",X"CD",X"8D",X"05",
		X"CD",X"BC",X"05",X"C9",X"DD",X"7E",X"00",X"3D",X"20",X"36",X"FD",X"7E",X"08",X"B7",X"20",X"06",
		X"3E",X"0F",X"CD",X"A9",X"08",X"C9",X"3D",X"4F",X"DD",X"7E",X"08",X"FD",X"86",X"09",X"DD",X"77",
		X"08",X"2A",X"02",X"10",X"06",X"00",X"09",X"09",X"46",X"23",X"66",X"68",X"23",X"23",X"BE",X"28",
		X"09",X"30",X"F9",X"CD",X"83",X"03",X"CD",X"A9",X"08",X"C9",X"23",X"7E",X"CD",X"A9",X"08",X"C9",
		X"DD",X"66",X"14",X"DD",X"6E",X"15",X"FD",X"56",X"02",X"FD",X"5E",X"01",X"AF",X"ED",X"52",X"38",
		X"0B",X"DD",X"75",X"15",X"7C",X"B7",X"28",X"04",X"CD",X"A9",X"08",X"C9",X"AF",X"DD",X"77",X"15",
		X"DD",X"77",X"00",X"CD",X"A9",X"08",X"AF",X"CD",X"C3",X"08",X"FD",X"35",X"18",X"C9",X"FD",X"7E",
		X"0A",X"B7",X"5F",X"20",X"0F",X"DD",X"7E",X"12",X"B7",X"C8",X"DD",X"6E",X"0F",X"DD",X"66",X"10",
		X"CD",X"04",X"09",X"C9",X"DD",X"7E",X"09",X"FD",X"86",X"0B",X"DD",X"77",X"09",X"4F",X"DD",X"7E",
		X"12",X"B7",X"C8",X"16",X"00",X"2A",X"04",X"10",X"1D",X"19",X"19",X"5E",X"23",X"66",X"6B",X"79",
		X"32",X"C9",X"81",X"11",X"05",X"00",X"19",X"BE",X"28",X"4D",X"30",X"FA",X"AF",X"32",X"CC",X"81",
		X"DD",X"E5",X"E5",X"DD",X"E1",X"DD",X"56",X"FF",X"DD",X"5E",X"FE",X"CB",X"7A",X"28",X"0C",X"7A",
		X"2F",X"57",X"7B",X"2F",X"5F",X"13",X"3E",X"01",X"32",X"CC",X"81",X"3A",X"C9",X"81",X"DD",X"96",
		X"FB",X"0E",X"00",X"CD",X"2D",X"04",X"EB",X"3A",X"CC",X"81",X"3D",X"20",X"06",X"21",X"00",X"00",
		X"ED",X"52",X"EB",X"DD",X"66",X"FD",X"DD",X"6E",X"FC",X"19",X"DD",X"E1",X"DD",X"5E",X"0F",X"DD",
		X"56",X"10",X"19",X"CD",X"04",X"09",X"C9",X"23",X"5E",X"23",X"66",X"6B",X"18",X"EE",X"FD",X"7E",
		X"0C",X"B7",X"C8",X"3D",X"4F",X"DD",X"7E",X"0A",X"FD",X"86",X"0D",X"DD",X"77",X"0A",X"06",X"00",
		X"2A",X"06",X"10",X"09",X"09",X"46",X"23",X"66",X"68",X"23",X"23",X"BE",X"28",X"09",X"30",X"F9",
		X"CD",X"83",X"03",X"CD",X"C3",X"08",X"C9",X"23",X"7E",X"CD",X"C3",X"08",X"C9",X"FD",X"7E",X"0E",
		X"B7",X"C8",X"3D",X"4F",X"DD",X"7E",X"0B",X"FD",X"86",X"0F",X"DD",X"77",X"0B",X"2A",X"08",X"10",
		X"06",X"00",X"09",X"09",X"46",X"23",X"66",X"68",X"23",X"23",X"BE",X"28",X"09",X"30",X"F9",X"CD",
		X"83",X"03",X"CD",X"82",X"09",X"C9",X"23",X"7E",X"CD",X"82",X"09",X"C9",X"FD",X"7E",X"12",X"FE",
		X"02",X"30",X"04",X"CD",X"44",X"09",X"C9",X"D6",X"02",X"4F",X"DD",X"7E",X"0D",X"FD",X"86",X"13",
		X"DD",X"77",X"0D",X"2A",X"0C",X"10",X"06",X"00",X"09",X"09",X"46",X"23",X"66",X"68",X"23",X"23",
		X"BE",X"28",X"08",X"30",X"F9",X"2B",X"7E",X"CD",X"44",X"09",X"C9",X"23",X"7E",X"CD",X"44",X"09",
		X"C9",X"FD",X"7E",X"10",X"FE",X"02",X"30",X"04",X"CD",X"92",X"09",X"C9",X"D6",X"02",X"4F",X"DD",
		X"7E",X"0C",X"FD",X"86",X"11",X"DD",X"77",X"0C",X"2A",X"0A",X"10",X"06",X"00",X"09",X"09",X"46",
		X"23",X"66",X"68",X"23",X"23",X"BE",X"28",X"08",X"30",X"F9",X"2B",X"7E",X"CD",X"92",X"09",X"C9",
		X"23",X"7E",X"CD",X"92",X"09",X"C9",X"DD",X"21",X"CE",X"06",X"AF",X"F5",X"DD",X"6E",X"00",X"DD",
		X"66",X"01",X"7C",X"B5",X"20",X"0A",X"F1",X"47",X"3A",X"C7",X"81",X"B0",X"32",X"C7",X"81",X"C9",
		X"DD",X"5E",X"04",X"DD",X"56",X"05",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"ED",X"B0",X"DD",X"6E",
		X"00",X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7A",X"B3",X"28",X"11",X"06",X"02",
		X"3E",X"00",X"77",X"BE",X"C2",X"C9",X"06",X"F6",X"FF",X"10",X"F7",X"23",X"1B",X"18",X"EB",X"DD",
		X"66",X"01",X"DD",X"6E",X"00",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7A",X"B3",X"28",X"06",X"36",
		X"00",X"23",X"1B",X"18",X"F6",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",
		X"03",X"7A",X"B3",X"28",X"14",X"7E",X"FE",X"00",X"20",X"2F",X"3E",X"01",X"77",X"BE",X"C2",X"C9",
		X"06",X"CB",X"27",X"30",X"F7",X"23",X"1B",X"18",X"E8",X"AF",X"DD",X"66",X"05",X"DD",X"6E",X"04",
		X"DD",X"56",X"01",X"DD",X"5E",X"00",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"ED",X"B0",X"47",X"F1",
		X"B0",X"11",X"07",X"00",X"DD",X"19",X"C3",X"2B",X"06",X"DD",X"7E",X"06",X"18",X"DC",X"00",X"80",
		X"00",X"02",X"00",X"80",X"10",X"00",X"82",X"00",X"02",X"00",X"80",X"10",X"00",X"00",X"DD",X"21",
		X"1A",X"07",X"16",X"00",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"DD",X"4E",X"00",X"DD",X"46",X"01",
		X"78",X"B1",X"28",X"1A",X"AF",X"86",X"23",X"0D",X"20",X"FB",X"05",X"20",X"F8",X"DD",X"BE",X"04",
		X"28",X"05",X"7A",X"DD",X"B6",X"05",X"57",X"01",X"06",X"00",X"DD",X"09",X"18",X"D6",X"7A",X"B7",
		X"C8",X"47",X"3A",X"C7",X"81",X"B0",X"32",X"C7",X"81",X"C9",X"00",X"10",X"00",X"00",X"8B",X"01",
		X"00",X"10",X"00",X"10",X"C9",X"02",X"00",X"10",X"00",X"20",X"D5",X"04",X"00",X"10",X"00",X"30",
		X"47",X"08",X"00",X"00",X"75",X"06",X"03",X"21",X"01",X"90",X"C5",X"E5",X"7E",X"B7",X"CA",X"E1",
		X"07",X"3D",X"CA",X"00",X"00",X"3D",X"20",X"05",X"18",X"11",X"C3",X"E1",X"07",X"3D",X"20",X"08",
		X"21",X"1F",X"80",X"CB",X"FE",X"C3",X"E1",X"07",X"3D",X"20",X"0A",X"21",X"1F",X"80",X"CB",X"BE",
		X"CD",X"BD",X"01",X"18",X"7C",X"3D",X"2A",X"00",X"10",X"07",X"CD",X"00",X"0B",X"7E",X"23",X"66",
		X"6F",X"E5",X"DD",X"E1",X"06",X"0A",X"21",X"43",X"80",X"11",X"19",X"00",X"7E",X"B7",X"20",X"5E",
		X"36",X"01",X"DD",X"7E",X"03",X"23",X"77",X"DD",X"7E",X"04",X"23",X"77",X"DD",X"7E",X"02",X"23",
		X"77",X"23",X"36",X"00",X"23",X"36",X"00",X"DD",X"7E",X"07",X"23",X"77",X"DD",X"7E",X"05",X"23",
		X"77",X"DD",X"7E",X"06",X"DD",X"E5",X"06",X"06",X"11",X"00",X"00",X"0E",X"00",X"07",X"30",X"0A",
		X"DD",X"56",X"08",X"DD",X"5E",X"09",X"DD",X"23",X"DD",X"23",X"23",X"72",X"23",X"73",X"10",X"E8",
		X"11",X"08",X"00",X"DD",X"19",X"DD",X"E5",X"D1",X"23",X"73",X"23",X"72",X"23",X"73",X"23",X"72",
		X"DD",X"E1",X"DD",X"66",X"01",X"DD",X"6E",X"00",X"7D",X"B4",X"20",X"95",X"18",X"03",X"19",X"10",
		X"9B",X"E1",X"23",X"C1",X"05",X"C2",X"3A",X"07",X"C9",X"D1",X"0F",X"EE",X"0E",X"18",X"0E",X"4D",
		X"0D",X"8E",X"0C",X"DA",X"0B",X"2F",X"0B",X"8F",X"0A",X"F7",X"09",X"68",X"09",X"E1",X"08",X"61",
		X"08",X"E9",X"07",X"77",X"07",X"0C",X"07",X"A7",X"06",X"47",X"06",X"ED",X"05",X"98",X"05",X"47",
		X"05",X"FB",X"04",X"B4",X"04",X"70",X"04",X"31",X"04",X"F4",X"03",X"BC",X"03",X"86",X"03",X"53",
		X"03",X"24",X"03",X"F6",X"02",X"CC",X"02",X"A4",X"02",X"7E",X"02",X"5A",X"02",X"38",X"02",X"18",
		X"02",X"FA",X"01",X"DE",X"01",X"C3",X"01",X"AA",X"01",X"92",X"01",X"7B",X"01",X"66",X"01",X"52",
		X"01",X"3F",X"01",X"2D",X"01",X"1C",X"01",X"0C",X"01",X"FD",X"00",X"EF",X"00",X"E1",X"00",X"D5",
		X"00",X"C9",X"00",X"BE",X"00",X"B3",X"00",X"A9",X"00",X"9F",X"00",X"96",X"00",X"8E",X"00",X"86",
		X"00",X"7F",X"00",X"77",X"00",X"71",X"00",X"6A",X"00",X"64",X"00",X"5F",X"00",X"59",X"00",X"54",
		X"00",X"50",X"00",X"4B",X"00",X"47",X"00",X"43",X"00",X"3F",X"00",X"3B",X"00",X"38",X"00",X"35",
		X"00",X"32",X"00",X"2F",X"00",X"2C",X"00",X"2A",X"00",X"27",X"00",X"26",X"00",X"24",X"00",X"22",
		X"00",X"20",X"00",X"1E",X"00",X"1C",X"00",X"1B",X"00",X"19",X"00",X"18",X"00",X"16",X"00",X"15",
		X"00",X"14",X"00",X"13",X"00",X"12",X"00",X"11",X"00",X"DD",X"BE",X"14",X"C8",X"DD",X"77",X"14",
		X"5F",X"21",X"08",X"80",X"DD",X"7E",X"01",X"FE",X"03",X"38",X"03",X"21",X"15",X"80",X"CD",X"00",
		X"0B",X"73",X"C9",X"DD",X"BE",X"16",X"C8",X"DD",X"77",X"16",X"16",X"00",X"21",X"EC",X"08",X"DD",
		X"5E",X"01",X"CB",X"23",X"CB",X"23",X"19",X"56",X"23",X"46",X"05",X"28",X"04",X"07",X"07",X"07",
		X"07",X"23",X"5E",X"23",X"66",X"6B",X"47",X"7E",X"A2",X"B0",X"77",X"C9",X"F0",X"01",X"0E",X"80",
		X"0F",X"02",X"0E",X"80",X"00",X"01",X"0F",X"80",X"F0",X"01",X"1E",X"80",X"0F",X"02",X"1E",X"80",
		X"00",X"01",X"1F",X"80",X"E5",X"6C",X"26",X"00",X"29",X"01",X"E9",X"07",X"09",X"4E",X"23",X"46",
		X"ED",X"43",X"CA",X"81",X"23",X"5E",X"23",X"56",X"60",X"69",X"AF",X"ED",X"52",X"5D",X"E1",X"65",
		X"CD",X"09",X"04",X"ED",X"5B",X"CA",X"81",X"6C",X"26",X"00",X"AF",X"EB",X"ED",X"52",X"EB",X"21",
		X"00",X"80",X"DD",X"7E",X"01",X"07",X"FE",X"06",X"38",X"03",X"21",X"0A",X"80",X"CD",X"00",X"0B",
		X"73",X"23",X"72",X"C9",X"DD",X"BE",X"13",X"C8",X"DD",X"77",X"13",X"16",X"00",X"21",X"6A",X"09",
		X"DD",X"5E",X"01",X"CB",X"23",X"CB",X"23",X"19",X"46",X"23",X"23",X"5E",X"23",X"66",X"6B",X"B7",
		X"78",X"20",X"03",X"B6",X"77",X"C9",X"2F",X"A6",X"77",X"C9",X"08",X"00",X"07",X"80",X"10",X"00",
		X"07",X"80",X"20",X"00",X"07",X"80",X"08",X"00",X"17",X"80",X"10",X"00",X"17",X"80",X"20",X"00",
		X"17",X"80",X"47",X"21",X"06",X"80",X"DD",X"7E",X"01",X"FE",X"03",X"38",X"03",X"21",X"16",X"80",
		X"70",X"C9",X"DD",X"BE",X"12",X"C8",X"DD",X"77",X"12",X"16",X"00",X"21",X"B8",X"09",X"DD",X"5E",
		X"01",X"CB",X"23",X"CB",X"23",X"19",X"46",X"23",X"23",X"5E",X"23",X"66",X"6B",X"B7",X"78",X"20",
		X"03",X"B6",X"77",X"C9",X"2F",X"A6",X"77",X"C9",X"01",X"00",X"07",X"80",X"02",X"00",X"07",X"80",
		X"04",X"00",X"07",X"80",X"01",X"00",X"17",X"80",X"02",X"00",X"17",X"80",X"04",X"00",X"17",X"80",
		X"21",X"00",X"80",X"11",X"01",X"80",X"36",X"00",X"01",X"F5",X"03",X"ED",X"B0",X"CD",X"BD",X"01",
		X"3A",X"00",X"90",X"E6",X"80",X"32",X"C8",X"81",X"C9",X"3A",X"00",X"90",X"B8",X"20",X"FA",X"3A",
		X"01",X"90",X"B8",X"20",X"F4",X"3A",X"02",X"90",X"B8",X"20",X"EE",X"3A",X"03",X"90",X"B8",X"20",
		X"E8",X"78",X"32",X"00",X"C0",X"C9",X"06",X"00",X"CD",X"7D",X"0A",X"0E",X"00",X"3E",X"AD",X"CD",
		X"66",X"0A",X"0E",X"01",X"3E",X"07",X"CD",X"66",X"0A",X"06",X"01",X"CD",X"7D",X"0A",X"0E",X"00",
		X"3E",X"AD",X"CD",X"66",X"0A",X"0E",X"01",X"3E",X"77",X"CD",X"66",X"0A",X"C9",X"CD",X"06",X"0A",
		X"16",X"10",X"3E",X"00",X"1E",X"FF",X"06",X"00",X"0E",X"00",X"CD",X"66",X"0A",X"2F",X"0E",X"01",
		X"CD",X"66",X"0A",X"06",X"01",X"32",X"80",X"0A",X"E6",X"7F",X"CD",X"66",X"0A",X"3A",X"80",X"0A",
		X"2F",X"0E",X"00",X"CD",X"66",X"0A",X"3C",X"E6",X"0F",X"47",X"07",X"07",X"07",X"07",X"B0",X"1D",
		X"20",X"FD",X"15",X"20",X"CF",X"C9",X"CD",X"7E",X"0A",X"32",X"7F",X"0A",X"AF",X"A9",X"28",X"09",
		X"36",X"0F",X"3A",X"7F",X"0A",X"DD",X"77",X"00",X"C9",X"36",X"0E",X"18",X"F5",X"C9",X"C9",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"85",X"6F",X"D0",X"24",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E0",X"34",X"C0",X"35",X"A7",X"36",X"D5",X"36",X"F3",X"36",X"01",X"37",X"09",X"37",X"00",X"00",
		X"00",X"55",X"00",X"00",X"08",X"0A",X"01",X"00",X"00",X"00",X"00",X"25",X"FF",X"05",X"F5",X"00",
		X"00",X"29",X"0A",X"05",X"E0",X"01",X"00",X"2C",X"1F",X"04",X"CB",X"02",X"00",X"31",X"34",X"03",
		X"BB",X"03",X"00",X"35",X"44",X"02",X"B5",X"04",X"00",X"38",X"45",X"01",X"00",X"FF",X"AE",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"48",X"0A",X"03",X"FF",X"01",X"7A",X"00",X"00",X"00",X"25",
		X"DD",X"00",X"0A",X"00",X"00",X"38",X"DD",X"00",X"0A",X"00",X"00",X"35",X"DD",X"00",X"64",X"00",
		X"00",X"31",X"DD",X"00",X"82",X"00",X"00",X"2C",X"DD",X"00",X"DC",X"00",X"00",X"35",X"DD",X"00",
		X"E6",X"00",X"00",X"38",X"DD",X"00",X"F0",X"00",X"00",X"25",X"DD",X"00",X"54",X"01",X"00",X"31",
		X"DD",X"00",X"5E",X"01",X"00",X"2C",X"DD",X"00",X"C2",X"01",X"00",X"25",X"DD",X"00",X"C2",X"01",
		X"00",X"35",X"DD",X"00",X"30",X"02",X"00",X"2C",X"DD",X"00",X"30",X"02",X"00",X"31",X"DD",X"00",
		X"94",X"02",X"00",X"25",X"DD",X"00",X"94",X"02",X"00",X"35",X"DD",X"00",X"02",X"03",X"00",X"2C",
		X"DD",X"00",X"02",X"03",X"00",X"31",X"DD",X"00",X"70",X"03",X"00",X"25",X"DD",X"00",X"70",X"03",
		X"00",X"35",X"DD",X"00",X"DE",X"03",X"00",X"2C",X"DD",X"00",X"DE",X"03",X"00",X"31",X"DD",X"00",
		X"42",X"04",X"00",X"25",X"DD",X"00",X"4C",X"04",X"00",X"35",X"DD",X"00",X"B0",X"04",X"00",X"31",
		X"DD",X"00",X"BA",X"04",X"00",X"2C",X"DD",X"00",X"1E",X"05",X"00",X"25",X"DD",X"00",X"1E",X"05",
		X"00",X"35",X"DD",X"00",X"8C",X"05",X"00",X"31",X"DD",X"00",X"96",X"05",X"00",X"2C",X"DD",X"00",
		X"FA",X"05",X"00",X"38",X"DD",X"00",X"FA",X"05",X"00",X"35",X"DD",X"00",X"04",X"06",X"00",X"25",
		X"DD",X"00",X"68",X"06",X"00",X"2C",X"DD",X"00",X"D6",X"06",X"00",X"35",X"DD",X"00",X"D6",X"06",
		X"00",X"38",X"DD",X"00",X"3A",X"07",X"00",X"31",X"DD",X"00",X"44",X"07",X"00",X"2C",X"DD",X"00",
		X"B2",X"07",X"00",X"25",X"DD",X"00",X"B2",X"07",X"00",X"35",X"DD",X"00",X"16",X"08",X"00",X"31",
		X"DD",X"00",X"20",X"08",X"00",X"2C",X"DD",X"00",X"84",X"08",X"00",X"25",X"DD",X"00",X"84",X"08",
		X"00",X"35",X"DD",X"00",X"F2",X"08",X"00",X"31",X"DD",X"00",X"06",X"09",X"00",X"2C",X"DD",X"00",
		X"60",X"09",X"00",X"25",X"DD",X"00",X"60",X"09",X"00",X"38",X"DD",X"00",X"6A",X"09",X"00",X"35",
		X"DD",X"00",X"CE",X"09",X"00",X"31",X"DD",X"00",X"D8",X"09",X"00",X"2C",X"DD",X"00",X"32",X"0A",
		X"00",X"35",X"DD",X"00",X"AA",X"0A",X"00",X"31",X"DD",X"00",X"B4",X"0A",X"00",X"2C",X"DD",X"00",
		X"0E",X"0B",X"00",X"38",X"DD",X"00",X"18",X"0B",X"00",X"25",X"DD",X"00",X"18",X"0B",X"00",X"35",
		X"DD",X"00",X"7C",X"0B",X"00",X"31",X"DD",X"00",X"90",X"0B",X"00",X"2C",X"DD",X"00",X"D6",X"0B",
		X"00",X"35",X"DD",X"00",X"58",X"0C",X"00",X"31",X"DD",X"00",X"6C",X"0C",X"00",X"2C",X"DD",X"00",
		X"A8",X"0C",X"00",X"38",X"DD",X"00",X"B2",X"0C",X"00",X"35",X"DD",X"00",X"C6",X"0C",X"00",X"25",
		X"DD",X"00",X"20",X"0D",X"00",X"31",X"DD",X"00",X"00",X"FF",X"70",X"0D",X"00",X"00",X"00",X"55",
		X"00",X"00",X"08",X"0D",X"01",X"7A",X"00",X"00",X"00",X"3A",X"1E",X"00",X"8A",X"00",X"00",X"36",
		X"2A",X"00",X"C0",X"00",X"00",X"33",X"24",X"00",X"92",X"01",X"00",X"31",X"4E",X"00",X"00",X"FF",
		X"06",X"03",X"00",X"00",X"01",X"89",X"00",X"00",X"08",X"09",X"01",X"00",X"00",X"00",X"00",X"2C",
		X"0C",X"00",X"18",X"00",X"00",X"2F",X"0C",X"00",X"30",X"00",X"00",X"34",X"0C",X"00",X"00",X"FF",
		X"D0",X"01",X"D0",X"13",X"02",X"6E",X"00",X"00",X"88",X"09",X"09",X"06",X"01",X"00",X"00",X"00",
		X"07",X"35",X"49",X"00",X"78",X"00",X"07",X"36",X"49",X"00",X"E8",X"00",X"07",X"38",X"49",X"00",
		X"68",X"01",X"07",X"3A",X"49",X"00",X"E0",X"03",X"07",X"3A",X"49",X"00",X"60",X"04",X"07",X"3C",
		X"49",X"00",X"E0",X"04",X"07",X"3D",X"49",X"00",X"50",X"05",X"07",X"3F",X"49",X"00",X"D0",X"05",
		X"07",X"3D",X"49",X"00",X"50",X"06",X"07",X"3D",X"49",X"00",X"C0",X"06",X"07",X"3C",X"49",X"00",
		X"48",X"07",X"07",X"3C",X"49",X"00",X"B8",X"07",X"07",X"3A",X"49",X"00",X"40",X"08",X"07",X"3A",
		X"49",X"00",X"A8",X"08",X"07",X"38",X"49",X"00",X"38",X"09",X"07",X"38",X"49",X"00",X"88",X"0B",
		X"07",X"35",X"49",X"00",X"10",X"0C",X"07",X"36",X"49",X"00",X"90",X"0C",X"07",X"38",X"49",X"00",
		X"10",X"0D",X"07",X"3A",X"49",X"00",X"A0",X"0F",X"07",X"3A",X"49",X"00",X"10",X"10",X"07",X"3C",
		X"49",X"00",X"80",X"10",X"07",X"3D",X"49",X"00",X"F8",X"10",X"07",X"3F",X"49",X"00",X"88",X"11",
		X"07",X"3D",X"49",X"00",X"00",X"12",X"07",X"3D",X"49",X"00",X"78",X"12",X"07",X"3C",X"49",X"00",
		X"00",X"13",X"07",X"3C",X"49",X"00",X"70",X"13",X"07",X"3A",X"49",X"00",X"F8",X"13",X"07",X"3A",
		X"49",X"00",X"60",X"14",X"07",X"38",X"49",X"00",X"D8",X"14",X"07",X"38",X"49",X"00",X"C8",X"15",
		X"07",X"41",X"49",X"00",X"48",X"16",X"07",X"41",X"49",X"00",X"50",X"17",X"07",X"41",X"49",X"00",
		X"B8",X"17",X"07",X"42",X"49",X"00",X"28",X"18",X"07",X"41",X"49",X"00",X"A8",X"18",X"07",X"41",
		X"49",X"00",X"18",X"19",X"07",X"3F",X"49",X"00",X"98",X"19",X"07",X"3F",X"49",X"00",X"E8",X"1A",
		X"07",X"3F",X"49",X"00",X"60",X"1B",X"07",X"41",X"49",X"00",X"D8",X"1B",X"07",X"42",X"49",X"00",
		X"60",X"1C",X"07",X"42",X"49",X"00",X"D0",X"1C",X"07",X"41",X"49",X"00",X"58",X"1D",X"07",X"41",
		X"49",X"00",X"D0",X"1E",X"07",X"41",X"49",X"00",X"48",X"1F",X"07",X"42",X"49",X"00",X"B0",X"1F",
		X"07",X"41",X"49",X"00",X"20",X"20",X"07",X"44",X"49",X"00",X"90",X"20",X"07",X"42",X"49",X"00",
		X"10",X"21",X"07",X"42",X"49",X"00",X"78",X"22",X"07",X"3F",X"49",X"00",X"F0",X"22",X"07",X"41",
		X"49",X"00",X"60",X"23",X"07",X"42",X"49",X"00",X"D0",X"23",X"07",X"42",X"49",X"00",X"40",X"24",
		X"07",X"41",X"49",X"00",X"C0",X"24",X"07",X"41",X"49",X"00",X"20",X"26",X"07",X"41",X"49",X"00",
		X"90",X"26",X"07",X"42",X"49",X"00",X"00",X"27",X"07",X"44",X"49",X"00",X"68",X"27",X"07",X"46",
		X"49",X"00",X"70",X"27",X"07",X"46",X"49",X"00",X"58",X"29",X"07",X"46",X"49",X"00",X"D0",X"29",
		X"07",X"44",X"49",X"00",X"70",X"2B",X"07",X"46",X"49",X"00",X"E8",X"2B",X"07",X"42",X"49",X"00",
		X"28",X"2C",X"07",X"3F",X"49",X"00",X"E0",X"2C",X"07",X"3D",X"49",X"00",X"00",X"FF",X"D0",X"31",
		X"F8",X"16",X"03",X"6E",X"00",X"00",X"88",X"09",X"09",X"06",X"01",X"00",X"77",X"00",X"00",X"19",
		X"49",X"00",X"77",X"00",X"00",X"23",X"49",X"00",X"77",X"00",X"00",X"25",X"49",X"00",X"5E",X"01",
		X"00",X"1E",X"49",X"00",X"E3",X"01",X"00",X"22",X"49",X"00",X"E3",X"01",X"00",X"25",X"49",X"00",
		X"6F",X"02",X"00",X"19",X"49",X"00",X"ED",X"02",X"00",X"22",X"49",X"00",X"ED",X"02",X"00",X"25",
		X"49",X"00",X"79",X"03",X"00",X"1E",X"49",X"00",X"F0",X"03",X"00",X"25",X"49",X"00",X"F7",X"03",
		X"00",X"22",X"49",X"00",X"67",X"04",X"00",X"19",X"49",X"00",X"DE",X"04",X"00",X"22",X"49",X"00",
		X"E5",X"04",X"00",X"25",X"49",X"00",X"63",X"05",X"00",X"1E",X"49",X"00",X"DA",X"05",X"00",X"24",
		X"49",X"00",X"DA",X"05",X"00",X"27",X"49",X"00",X"58",X"06",X"00",X"1B",X"49",X"00",X"C8",X"06",
		X"00",X"24",X"49",X"00",X"C8",X"06",X"00",X"27",X"49",X"00",X"46",X"07",X"00",X"20",X"49",X"00",
		X"C4",X"07",X"00",X"24",X"49",X"00",X"C4",X"07",X"00",X"27",X"49",X"00",X"34",X"08",X"00",X"1B",
		X"49",X"00",X"B2",X"08",X"00",X"27",X"49",X"00",X"B9",X"08",X"00",X"24",X"49",X"00",X"29",X"09",
		X"00",X"1D",X"49",X"00",X"A0",X"09",X"00",X"20",X"49",X"00",X"A0",X"09",X"00",X"25",X"49",X"00",
		X"25",X"0A",X"00",X"19",X"49",X"00",X"9C",X"0A",X"00",X"20",X"49",X"00",X"9C",X"0A",X"00",X"25",
		X"49",X"00",X"1A",X"0B",X"00",X"1D",X"49",X"00",X"08",X"0C",X"00",X"19",X"49",X"00",X"08",X"0C",
		X"00",X"23",X"49",X"00",X"08",X"0C",X"00",X"25",X"49",X"00",X"12",X"0D",X"00",X"1E",X"49",X"00",
		X"89",X"0D",X"00",X"22",X"49",X"00",X"89",X"0D",X"00",X"25",X"49",X"00",X"0E",X"0E",X"00",X"19",
		X"49",X"00",X"8C",X"0E",X"00",X"22",X"49",X"00",X"8C",X"0E",X"00",X"25",X"49",X"00",X"11",X"0F",
		X"00",X"1E",X"49",X"00",X"88",X"0F",X"00",X"22",X"49",X"00",X"88",X"0F",X"00",X"25",X"49",X"00",
		X"1B",X"10",X"00",X"19",X"49",X"00",X"92",X"10",X"00",X"22",X"49",X"00",X"92",X"10",X"00",X"25",
		X"49",X"00",X"17",X"11",X"00",X"1E",X"49",X"00",X"79",X"11",X"00",X"24",X"49",X"00",X"80",X"11",
		X"00",X"27",X"49",X"00",X"05",X"12",X"00",X"1B",X"49",X"00",X"75",X"12",X"00",X"24",X"49",X"00",
		X"75",X"12",X"00",X"27",X"49",X"00",X"FA",X"12",X"00",X"20",X"49",X"00",X"6A",X"13",X"00",X"24",
		X"49",X"00",X"6A",X"13",X"00",X"27",X"49",X"00",X"EF",X"13",X"00",X"1B",X"49",X"00",X"58",X"14",
		X"00",X"27",X"49",X"00",X"66",X"14",X"00",X"24",X"49",X"00",X"DD",X"14",X"00",X"1D",X"49",X"00",
		X"54",X"15",X"00",X"20",X"49",X"00",X"5B",X"15",X"00",X"25",X"49",X"00",X"D9",X"15",X"00",X"19",
		X"49",X"00",X"49",X"16",X"00",X"25",X"49",X"00",X"50",X"16",X"00",X"20",X"49",X"00",X"C7",X"16",
		X"00",X"1D",X"49",X"00",X"45",X"17",X"00",X"20",X"49",X"00",X"45",X"17",X"00",X"25",X"49",X"00",
		X"C3",X"17",X"00",X"19",X"49",X"00",X"33",X"18",X"00",X"20",X"49",X"00",X"33",X"18",X"00",X"25",
		X"49",X"00",X"AA",X"18",X"00",X"1E",X"49",X"00",X"2F",X"19",X"00",X"23",X"49",X"00",X"2F",X"19",
		X"00",X"27",X"49",X"00",X"A6",X"19",X"00",X"1B",X"49",X"00",X"16",X"1A",X"00",X"23",X"49",X"00",
		X"1D",X"1A",X"00",X"27",X"49",X"00",X"55",X"1A",X"00",X"23",X"49",X"00",X"94",X"1A",X"00",X"1E",
		X"49",X"00",X"0B",X"1B",X"00",X"23",X"49",X"00",X"0B",X"1B",X"00",X"27",X"49",X"00",X"7B",X"1B",
		X"00",X"1B",X"49",X"00",X"E4",X"1B",X"00",X"23",X"49",X"00",X"F2",X"1B",X"00",X"27",X"49",X"00",
		X"70",X"1C",X"00",X"20",X"49",X"00",X"D9",X"1C",X"00",X"25",X"49",X"00",X"E0",X"1C",X"00",X"29",
		X"49",X"00",X"49",X"1D",X"00",X"1D",X"49",X"00",X"C7",X"1D",X"00",X"25",X"49",X"00",X"C7",X"1D",
		X"00",X"29",X"49",X"00",X"3E",X"1E",X"00",X"20",X"49",X"00",X"C3",X"1E",X"00",X"25",X"49",X"00",
		X"C3",X"1E",X"00",X"29",X"49",X"00",X"41",X"1F",X"00",X"1D",X"49",X"00",X"B8",X"1F",X"00",X"25",
		X"49",X"00",X"BF",X"1F",X"00",X"29",X"49",X"00",X"28",X"20",X"00",X"1E",X"49",X"00",X"9F",X"20",
		X"00",X"23",X"49",X"00",X"9F",X"20",X"00",X"27",X"49",X"00",X"16",X"21",X"00",X"1B",X"49",X"00",
		X"8D",X"21",X"00",X"23",X"49",X"00",X"94",X"21",X"00",X"27",X"49",X"00",X"04",X"22",X"00",X"1E",
		X"49",X"00",X"74",X"22",X"00",X"23",X"49",X"00",X"7B",X"22",X"00",X"27",X"49",X"00",X"EB",X"22",
		X"00",X"1B",X"49",X"00",X"5B",X"23",X"00",X"23",X"49",X"00",X"5B",X"23",X"00",X"27",X"49",X"00",
		X"D2",X"23",X"00",X"20",X"49",X"00",X"49",X"24",X"00",X"25",X"49",X"00",X"57",X"24",X"00",X"29",
		X"49",X"00",X"B9",X"24",X"00",X"1D",X"49",X"00",X"30",X"25",X"00",X"25",X"49",X"00",X"37",X"25",
		X"00",X"29",X"49",X"00",X"A0",X"25",X"00",X"20",X"49",X"00",X"17",X"26",X"00",X"25",X"49",X"00",
		X"1E",X"26",X"00",X"29",X"49",X"00",X"95",X"26",X"00",X"1D",X"49",X"00",X"FE",X"26",X"00",X"25",
		X"49",X"00",X"FE",X"26",X"00",X"29",X"49",X"00",X"91",X"27",X"00",X"1E",X"49",X"00",X"91",X"27",
		X"00",X"22",X"49",X"00",X"98",X"27",X"00",X"25",X"49",X"00",X"4A",X"29",X"00",X"20",X"49",X"00",
		X"4A",X"29",X"00",X"24",X"49",X"00",X"4A",X"29",X"00",X"27",X"49",X"00",X"3B",X"2B",X"00",X"22",
		X"49",X"00",X"D5",X"2B",X"00",X"1E",X"49",X"00",X"0D",X"2C",X"00",X"1B",X"49",X"00",X"D8",X"2C",
		X"00",X"19",X"49",X"00",X"00",X"FF",X"80",X"2D",X"00",X"00",X"03",X"6E",X"00",X"00",X"88",X"09",
		X"09",X"06",X"01",X"00",X"81",X"01",X"00",X"12",X"49",X"00",X"6F",X"02",X"00",X"0D",X"49",X"00",
		X"79",X"03",X"00",X"12",X"49",X"00",X"67",X"04",X"00",X"0D",X"49",X"00",X"63",X"05",X"00",X"12",
		X"49",X"00",X"3C",X"06",X"00",X"0F",X"49",X"00",X"38",X"07",X"00",X"14",X"49",X"00",X"3B",X"08",
		X"00",X"0F",X"49",X"00",X"22",X"09",X"00",X"11",X"49",X"00",X"25",X"0A",X"00",X"0D",X"49",X"00",
		X"1A",X"0B",X"00",X"11",X"49",X"00",X"20",X"0D",X"00",X"12",X"49",X"00",X"23",X"0E",X"00",X"0D",
		X"49",X"00",X"1F",X"0F",X"00",X"12",X"49",X"00",X"1B",X"10",X"00",X"0D",X"49",X"00",X"09",X"11",
		X"00",X"12",X"49",X"00",X"FE",X"11",X"00",X"0F",X"49",X"00",X"08",X"13",X"00",X"14",X"49",X"00",
		X"FD",X"13",X"00",X"0F",X"49",X"00",X"EB",X"14",X"00",X"11",X"49",X"00",X"EE",X"15",X"00",X"0D",
		X"49",X"00",X"E3",X"16",X"00",X"11",X"49",X"00",X"BC",X"17",X"00",X"0D",X"49",X"00",X"B1",X"18",
		X"00",X"12",X"49",X"00",X"A6",X"19",X"00",X"0F",X"49",X"00",X"9B",X"1A",X"00",X"12",X"49",X"00",
		X"74",X"1B",X"00",X"0F",X"49",X"00",X"5B",X"1C",X"00",X"11",X"49",X"00",X"5E",X"1D",X"00",X"0D",
		X"49",X"00",X"61",X"1E",X"00",X"11",X"49",X"00",X"4F",X"1F",X"00",X"0D",X"49",X"00",X"2F",X"20",
		X"00",X"12",X"49",X"00",X"1D",X"21",X"00",X"0F",X"49",X"00",X"0B",X"22",X"00",X"12",X"49",X"00",
		X"F2",X"22",X"00",X"0F",X"49",X"00",X"D9",X"23",X"00",X"11",X"49",X"00",X"B9",X"24",X"00",X"0D",
		X"49",X"00",X"B5",X"25",X"00",X"11",X"49",X"00",X"9C",X"26",X"00",X"0D",X"49",X"00",X"8A",X"27",
		X"00",X"12",X"49",X"00",X"7B",X"29",X"00",X"14",X"49",X"00",X"00",X"FF",X"59",X"2E",X"00",X"00",
		X"14",X"3A",X"00",X"FF",X"88",X"0C",X"04",X"00",X"01",X"00",X"00",X"00",X"00",X"2A",X"49",X"00",
		X"6C",X"00",X"00",X"2C",X"49",X"00",X"BA",X"00",X"00",X"1E",X"49",X"00",X"BA",X"00",X"00",X"2E",
		X"49",X"00",X"5C",X"01",X"00",X"22",X"49",X"00",X"5C",X"01",X"00",X"25",X"49",X"00",X"62",X"01",
		X"00",X"31",X"49",X"00",X"0A",X"02",X"00",X"19",X"49",X"00",X"0A",X"02",X"00",X"31",X"49",X"00",
		X"AC",X"02",X"00",X"22",X"49",X"00",X"AC",X"02",X"00",X"33",X"49",X"00",X"B2",X"02",X"00",X"25",
		X"49",X"00",X"54",X"03",X"00",X"1E",X"49",X"00",X"54",X"03",X"00",X"31",X"49",X"00",X"F6",X"03",
		X"00",X"22",X"49",X"00",X"F6",X"03",X"00",X"25",X"49",X"00",X"FC",X"03",X"00",X"2E",X"49",X"00",
		X"9E",X"04",X"00",X"19",X"49",X"00",X"A4",X"04",X"00",X"2A",X"49",X"00",X"46",X"05",X"00",X"22",
		X"49",X"00",X"46",X"05",X"00",X"25",X"49",X"00",X"46",X"05",X"00",X"2C",X"49",X"00",X"E8",X"05",
		X"00",X"1E",X"49",X"00",X"F4",X"05",X"00",X"2E",X"49",X"00",X"90",X"06",X"00",X"22",X"49",X"00",
		X"96",X"06",X"00",X"25",X"49",X"00",X"96",X"06",X"00",X"2E",X"49",X"00",X"26",X"07",X"00",X"19",
		X"49",X"00",X"38",X"07",X"00",X"2C",X"49",X"00",X"D4",X"07",X"00",X"22",X"49",X"00",X"D4",X"07",
		X"00",X"25",X"49",X"00",X"D4",X"07",X"00",X"2A",X"49",X"00",X"82",X"08",X"00",X"1D",X"49",X"00",
		X"88",X"08",X"00",X"2C",X"49",X"00",X"2A",X"09",X"00",X"25",X"49",X"00",X"30",X"09",X"00",X"20",
		X"49",X"00",X"D8",X"09",X"00",X"19",X"49",X"00",X"68",X"0A",X"00",X"25",X"49",X"00",X"6E",X"0A",
		X"00",X"20",X"49",X"00",X"6E",X"0A",X"00",X"2A",X"49",X"00",X"DA",X"0A",X"00",X"2C",X"49",X"00",
		X"1C",X"0B",X"00",X"2E",X"49",X"00",X"22",X"0B",X"00",X"1E",X"49",X"00",X"BE",X"0B",X"00",X"22",
		X"49",X"00",X"BE",X"0B",X"00",X"25",X"49",X"00",X"C4",X"0B",X"00",X"31",X"49",X"00",X"6C",X"0C",
		X"00",X"19",X"49",X"00",X"6C",X"0C",X"00",X"31",X"49",X"00",X"0E",X"0D",X"00",X"22",X"49",X"00",
		X"0E",X"0D",X"00",X"25",X"49",X"00",X"6E",X"0D",X"00",X"33",X"49",X"00",X"AA",X"0D",X"00",X"1E",
		X"49",X"00",X"AA",X"0D",X"00",X"31",X"49",X"00",X"40",X"0E",X"00",X"22",X"49",X"00",X"40",X"0E",
		X"00",X"25",X"49",X"00",X"46",X"0E",X"00",X"2E",X"49",X"00",X"E2",X"0E",X"00",X"19",X"49",X"00",
		X"EE",X"0E",X"00",X"2A",X"49",X"00",X"8A",X"0F",X"00",X"22",X"49",X"00",X"8A",X"0F",X"00",X"25",
		X"49",X"00",X"90",X"0F",X"00",X"2C",X"49",X"00",X"38",X"10",X"00",X"2E",X"49",X"00",X"44",X"10",
		X"00",X"1E",X"49",X"00",X"DA",X"10",X"00",X"24",X"49",X"00",X"DA",X"10",X"00",X"27",X"49",X"00",
		X"E0",X"10",X"00",X"2E",X"49",X"00",X"82",X"11",X"00",X"1B",X"49",X"00",X"88",X"11",X"00",X"2C",
		X"49",X"00",X"42",X"12",X"00",X"20",X"49",X"00",X"4E",X"12",X"00",X"2C",X"49",X"00",X"54",X"12",
		X"00",X"25",X"49",X"00",X"EA",X"12",X"00",X"1E",X"49",X"00",X"F0",X"12",X"00",X"2A",X"49",X"00",
		X"8C",X"13",X"00",X"22",X"49",X"00",X"8C",X"13",X"00",X"25",X"49",X"00",X"40",X"14",X"00",X"19",
		X"49",X"00",X"D6",X"14",X"00",X"22",X"49",X"00",X"DC",X"14",X"00",X"25",X"49",X"00",X"DC",X"14",
		X"00",X"2A",X"49",X"00",X"42",X"15",X"00",X"2C",X"49",X"00",X"78",X"15",X"00",X"2E",X"49",X"00",
		X"7E",X"15",X"00",X"1E",X"49",X"00",X"1A",X"16",X"00",X"22",X"49",X"00",X"1A",X"16",X"00",X"25",
		X"49",X"00",X"1A",X"16",X"00",X"31",X"49",X"00",X"BC",X"16",X"00",X"19",X"49",X"00",X"C2",X"16",
		X"00",X"31",X"49",X"00",X"5E",X"17",X"00",X"22",X"49",X"00",X"5E",X"17",X"00",X"25",X"49",X"00",
		X"BE",X"17",X"00",X"33",X"49",X"00",X"FA",X"17",X"00",X"1E",X"49",X"00",X"FA",X"17",X"00",X"31",
		X"49",X"00",X"96",X"18",X"00",X"25",X"49",X"00",X"9C",X"18",X"00",X"22",X"49",X"00",X"9C",X"18",
		X"00",X"2E",X"49",X"00",X"32",X"19",X"00",X"19",X"49",X"00",X"3E",X"19",X"00",X"2A",X"49",X"00",
		X"DA",X"19",X"00",X"22",X"49",X"00",X"DA",X"19",X"00",X"25",X"49",X"00",X"DA",X"19",X"00",X"2C",
		X"49",X"00",X"82",X"1A",X"00",X"1E",X"49",X"00",X"88",X"1A",X"00",X"2E",X"49",X"00",X"1E",X"1B",
		X"00",X"24",X"49",X"00",X"1E",X"1B",X"00",X"27",X"49",X"00",X"24",X"1B",X"00",X"2E",X"49",X"00",
		X"C0",X"1B",X"00",X"1B",X"49",X"00",X"CC",X"1B",X"00",X"2C",X"49",X"00",X"62",X"1C",X"00",X"24",
		X"49",X"00",X"62",X"1C",X"00",X"27",X"49",X"00",X"68",X"1C",X"00",X"2A",X"49",X"00",X"04",X"1D",
		X"00",X"1D",X"49",X"00",X"04",X"1D",X"00",X"2C",X"49",X"00",X"A6",X"1D",X"00",X"20",X"49",X"00",
		X"A6",X"1D",X"00",X"25",X"49",X"00",X"48",X"1E",X"00",X"19",X"49",X"00",X"D8",X"1E",X"00",X"20",
		X"49",X"00",X"D8",X"1E",X"00",X"25",X"49",X"00",X"DE",X"1E",X"00",X"2A",X"49",X"00",X"38",X"1F",
		X"00",X"2C",X"49",X"00",X"80",X"1F",X"00",X"1E",X"49",X"00",X"86",X"1F",X"00",X"2E",X"49",X"00",
		X"2E",X"20",X"00",X"22",X"49",X"00",X"2E",X"20",X"00",X"25",X"49",X"00",X"2E",X"20",X"00",X"31",
		X"49",X"00",X"CA",X"20",X"00",X"19",X"49",X"00",X"D6",X"20",X"00",X"31",X"49",X"00",X"6C",X"21",
		X"00",X"22",X"49",X"00",X"6C",X"21",X"00",X"25",X"49",X"00",X"D2",X"21",X"00",X"33",X"49",X"00",
		X"0E",X"22",X"00",X"1E",X"49",X"00",X"0E",X"22",X"00",X"31",X"49",X"00",X"B0",X"22",X"00",X"22",
		X"49",X"00",X"B0",X"22",X"00",X"25",X"49",X"00",X"B0",X"22",X"00",X"2E",X"49",X"00",X"4C",X"23",
		X"00",X"19",X"49",X"00",X"58",X"23",X"00",X"2A",X"49",X"00",X"F4",X"23",X"00",X"22",X"49",X"00",
		X"F4",X"23",X"00",X"25",X"49",X"00",X"F4",X"23",X"00",X"2C",X"49",X"00",X"96",X"24",X"00",X"1D",
		X"49",X"00",X"9C",X"24",X"00",X"2E",X"49",X"00",X"32",X"25",X"00",X"20",X"49",X"00",X"32",X"25",
		X"00",X"25",X"49",X"00",X"38",X"25",X"00",X"2E",X"49",X"00",X"CE",X"25",X"00",X"19",X"49",X"00",
		X"DA",X"25",X"00",X"2C",X"49",X"00",X"76",X"26",X"00",X"20",X"49",X"00",X"76",X"26",X"00",X"25",
		X"49",X"00",X"76",X"26",X"00",X"2C",X"49",X"00",X"0C",X"27",X"00",X"1E",X"49",X"00",X"18",X"27",
		X"00",X"2A",X"49",X"00",X"AE",X"27",X"00",X"22",X"49",X"00",X"AE",X"27",X"00",X"25",X"49",X"00",
		X"56",X"28",X"00",X"19",X"49",X"00",X"F2",X"28",X"00",X"22",X"49",X"00",X"F2",X"28",X"00",X"25",
		X"49",X"00",X"94",X"29",X"00",X"1E",X"49",X"00",X"A0",X"29",X"00",X"33",X"49",X"00",X"30",X"2A",
		X"00",X"23",X"49",X"00",X"36",X"2A",X"00",X"27",X"49",X"00",X"CC",X"2A",X"00",X"1B",X"49",X"00",
		X"D2",X"2A",X"00",X"33",X"49",X"00",X"6E",X"2B",X"00",X"23",X"49",X"00",X"74",X"2B",X"00",X"27",
		X"49",X"00",X"0A",X"2C",X"00",X"1E",X"49",X"00",X"16",X"2C",X"00",X"36",X"49",X"00",X"A6",X"2C",
		X"00",X"23",X"49",X"00",X"A6",X"2C",X"00",X"27",X"49",X"00",X"AC",X"2C",X"00",X"36",X"49",X"00",
		X"42",X"2D",X"00",X"1B",X"49",X"00",X"D2",X"2D",X"00",X"23",X"49",X"00",X"D2",X"2D",X"00",X"27",
		X"49",X"00",X"D8",X"2D",X"00",X"33",X"49",X"00",X"68",X"2E",X"00",X"1E",X"49",X"00",X"74",X"2E",
		X"00",X"31",X"49",X"00",X"0A",X"2F",X"00",X"22",X"49",X"00",X"0A",X"2F",X"00",X"25",X"49",X"00",
		X"10",X"2F",X"00",X"31",X"49",X"00",X"B8",X"2F",X"00",X"19",X"49",X"00",X"BE",X"2F",X"00",X"2E",
		X"49",X"00",X"4E",X"30",X"00",X"25",X"49",X"00",X"54",X"30",X"00",X"22",X"49",X"00",X"5A",X"30",
		X"00",X"2A",X"49",X"00",X"FC",X"30",X"00",X"1D",X"49",X"00",X"FC",X"30",X"00",X"2C",X"49",X"00",
		X"8C",X"31",X"00",X"20",X"49",X"00",X"8C",X"31",X"00",X"25",X"49",X"00",X"2E",X"32",X"00",X"19",
		X"49",X"00",X"C4",X"32",X"00",X"25",X"49",X"00",X"C4",X"32",X"00",X"2A",X"49",X"00",X"CA",X"32",
		X"00",X"20",X"49",X"00",X"2A",X"33",X"00",X"2C",X"49",X"00",X"6C",X"33",X"00",X"1E",X"49",X"00",
		X"6C",X"33",X"00",X"2E",X"49",X"00",X"FC",X"33",X"00",X"22",X"49",X"00",X"02",X"34",X"00",X"25",
		X"49",X"00",X"08",X"34",X"00",X"31",X"49",X"00",X"9E",X"34",X"00",X"19",X"49",X"00",X"A4",X"34",
		X"00",X"31",X"49",X"00",X"34",X"35",X"00",X"22",X"49",X"00",X"34",X"35",X"00",X"25",X"49",X"00",
		X"9A",X"35",X"00",X"33",X"49",X"00",X"D6",X"35",X"00",X"1E",X"49",X"00",X"D6",X"35",X"00",X"31",
		X"49",X"00",X"66",X"36",X"00",X"22",X"49",X"00",X"66",X"36",X"00",X"25",X"49",X"00",X"6C",X"36",
		X"00",X"2E",X"49",X"00",X"F6",X"36",X"00",X"19",X"49",X"00",X"08",X"37",X"00",X"2A",X"49",X"00",
		X"98",X"37",X"00",X"22",X"49",X"00",X"9E",X"37",X"00",X"25",X"49",X"00",X"A4",X"37",X"00",X"2C",
		X"49",X"00",X"2E",X"38",X"00",X"1E",X"49",X"00",X"3A",X"38",X"00",X"2E",X"49",X"00",X"D0",X"38",
		X"00",X"24",X"49",X"00",X"D0",X"38",X"00",X"27",X"49",X"00",X"DC",X"38",X"00",X"2E",X"49",X"00",
		X"60",X"39",X"00",X"1D",X"49",X"00",X"72",X"39",X"00",X"2C",X"49",X"00",X"02",X"3A",X"00",X"20",
		X"49",X"00",X"02",X"3A",X"00",X"25",X"49",X"00",X"08",X"3A",X"00",X"2C",X"49",X"00",X"9E",X"3A",
		X"00",X"1E",X"49",X"00",X"A4",X"3A",X"00",X"2A",X"49",X"00",X"3A",X"3B",X"00",X"22",X"49",X"00",
		X"3A",X"3B",X"00",X"25",X"49",X"00",X"E2",X"3B",X"00",X"19",X"49",X"00",X"00",X"FF",X"96",X"3C",
		X"00",X"00",X"04",X"00",X"00",X"00",X"D8",X"0A",X"08",X"13",X"03",X"E9",X"02",X"F7",X"01",X"00",
		X"00",X"00",X"00",X"35",X"61",X"00",X"00",X"FF",X"C6",X"02",X"00",X"00",X"04",X"00",X"00",X"00",
		X"D8",X"0A",X"08",X"13",X"03",X"E9",X"02",X"F7",X"01",X"00",X"00",X"00",X"00",X"2C",X"61",X"00",
		X"00",X"FF",X"DA",X"02",X"00",X"00",X"0D",X"DF",X"02",X"00",X"48",X"0A",X"03",X"8B",X"01",X"3E",
		X"00",X"00",X"00",X"33",X"25",X"00",X"00",X"FF",X"B2",X"02",X"00",X"00",X"0D",X"DF",X"02",X"00",
		X"48",X"0A",X"03",X"8B",X"01",X"3E",X"00",X"00",X"00",X"31",X"25",X"00",X"00",X"FF",X"8A",X"02",
		X"00",X"00",X"03",X"00",X"00",X"00",X"68",X"0B",X"06",X"12",X"03",X"57",X"01",X"46",X"00",X"00",
		X"00",X"2F",X"96",X"00",X"00",X"FF",X"B5",X"02",X"00",X"00",X"04",X"00",X"00",X"00",X"B4",X"0A",
		X"01",X"15",X"02",X"0D",X"02",X"10",X"01",X"00",X"00",X"00",X"00",X"20",X"AA",X"00",X"00",X"FF",
		X"08",X"02",X"00",X"00",X"02",X"80",X"00",X"00",X"08",X"4B",X"01",X"00",X"00",X"00",X"00",X"31",
		X"32",X"00",X"64",X"00",X"00",X"36",X"28",X"00",X"CD",X"00",X"00",X"3A",X"28",X"00",X"3B",X"01",
		X"00",X"3D",X"32",X"00",X"9F",X"01",X"00",X"3A",X"28",X"00",X"08",X"02",X"00",X"36",X"23",X"00",
		X"76",X"02",X"00",X"31",X"37",X"00",X"DF",X"02",X"00",X"36",X"23",X"00",X"3E",X"03",X"00",X"3A",
		X"2D",X"00",X"A2",X"03",X"00",X"3D",X"23",X"00",X"00",X"FF",X"37",X"05",X"00",X"00",X"01",X"00",
		X"00",X"00",X"E8",X"06",X"05",X"03",X"05",X"03",X"03",X"25",X"01",X"42",X"00",X"00",X"BA",X"29",
		X"90",X"01",X"00",X"00",X"44",X"40",X"90",X"01",X"00",X"FF",X"08",X"04",X"00",X"00",X"04",X"00",
		X"00",X"00",X"48",X"06",X"02",X"FD",X"02",X"47",X"00",X"00",X"00",X"1D",X"5F",X"01",X"00",X"FF",
		X"1C",X"02",X"00",X"00",X"03",X"5A",X"00",X"00",X"08",X"0A",X"01",X"00",X"00",X"00",X"9E",X"4E",
		X"0A",X"00",X"23",X"00",X"D2",X"4C",X"0A",X"00",X"46",X"00",X"9E",X"4E",X"0A",X"00",X"69",X"00",
		X"D2",X"4C",X"0A",X"00",X"85",X"00",X"9E",X"4E",X"0A",X"00",X"00",X"FF",X"B2",X"01",X"00",X"00",
		X"04",X"00",X"00",X"00",X"94",X"0A",X"05",X"21",X"01",X"8B",X"01",X"00",X"00",X"00",X"00",X"2E",
		X"1F",X"00",X"00",X"FF",X"7A",X"03",X"D4",X"1E",X"04",X"74",X"00",X"00",X"58",X"0A",X"02",X"02",
		X"03",X"0A",X"01",X"00",X"00",X"00",X"00",X"23",X"EC",X"03",X"00",X"00",X"00",X"24",X"EC",X"03",
		X"00",X"FF",X"1A",X"09",X"00",X"00",X"04",X"5F",X"00",X"00",X"C8",X"0A",X"0A",X"1A",X"06",X"FF",
		X"01",X"00",X"00",X"00",X"00",X"16",X"0F",X"04",X"1E",X"00",X"00",X"20",X"0F",X"04",X"1E",X"00",
		X"00",X"27",X"0F",X"04",X"28",X"00",X"00",X"29",X"0F",X"04",X"32",X"00",X"00",X"19",X"0F",X"04",
		X"3C",X"00",X"00",X"1B",X"0F",X"04",X"00",X"FF",X"08",X"07",X"6C",X"1F",X"03",X"9E",X"00",X"00",
		X"B4",X"0A",X"09",X"00",X"02",X"16",X"03",X"0A",X"01",X"00",X"00",X"00",X"C0",X"45",X"0B",X"00",
		X"0A",X"00",X"E0",X"41",X"0B",X"00",X"46",X"00",X"40",X"55",X"0B",X"00",X"46",X"00",X"00",X"5D",
		X"0B",X"00",X"50",X"00",X"80",X"4D",X"0B",X"00",X"78",X"00",X"C0",X"45",X"0B",X"00",X"96",X"00",
		X"A0",X"49",X"0B",X"00",X"AA",X"00",X"40",X"55",X"0B",X"00",X"DC",X"00",X"A0",X"49",X"0B",X"00",
		X"36",X"01",X"20",X"59",X"0B",X"00",X"40",X"01",X"00",X"3E",X"0B",X"00",X"FE",X"01",X"40",X"36",
		X"0B",X"00",X"A8",X"02",X"00",X"3E",X"0B",X"00",X"00",X"FF",X"3E",X"08",X"A6",X"1F",X"03",X"74",
		X"00",X"00",X"14",X"0A",X"04",X"0A",X"01",X"00",X"00",X"00",X"00",X"1E",X"78",X"00",X"14",X"00",
		X"00",X"24",X"78",X"00",X"BE",X"00",X"00",X"25",X"50",X"00",X"04",X"01",X"00",X"24",X"64",X"00",
		X"40",X"01",X"00",X"1D",X"46",X"00",X"68",X"01",X"00",X"1B",X"78",X"00",X"CC",X"01",X"00",X"22",
		X"46",X"00",X"00",X"FF",X"FA",X"0A",X"0A",X"20",X"03",X"9E",X"00",X"00",X"84",X"0A",X"09",X"00",
		X"01",X"00",X"00",X"00",X"80",X"0F",X"0B",X"00",X"0A",X"00",X"00",X"00",X"0B",X"00",X"14",X"00",
		X"20",X"1B",X"0B",X"00",X"1E",X"00",X"E0",X"03",X"0B",X"00",X"1E",X"00",X"A0",X"0B",X"0B",X"00",
		X"28",X"00",X"00",X"00",X"0B",X"00",X"5A",X"00",X"A0",X"0B",X"0B",X"00",X"64",X"00",X"80",X"2E",
		X"0B",X"00",X"8C",X"00",X"80",X"0F",X"0B",X"00",X"96",X"00",X"60",X"13",X"0B",X"00",X"AA",X"00",
		X"00",X"00",X"0B",X"00",X"D2",X"00",X"C0",X"26",X"0B",X"00",X"FA",X"00",X"40",X"17",X"0B",X"00",
		X"04",X"01",X"60",X"13",X"0B",X"00",X"00",X"FF",X"0C",X"08",X"00",X"00",X"03",X"74",X"00",X"00",
		X"98",X"0A",X"09",X"00",X"04",X"0A",X"01",X"00",X"00",X"00",X"95",X"4A",X"32",X"00",X"00",X"00",
		X"6A",X"55",X"50",X"00",X"14",X"00",X"95",X"57",X"0A",X"00",X"32",X"00",X"BF",X"59",X"64",X"00",
		X"64",X"00",X"95",X"57",X"6E",X"00",X"AA",X"00",X"6A",X"55",X"78",X"00",X"DC",X"00",X"BF",X"59",
		X"0A",X"00",X"E6",X"00",X"BF",X"59",X"5A",X"00",X"04",X"01",X"95",X"57",X"78",X"00",X"5E",X"01",
		X"6A",X"55",X"96",X"00",X"A4",X"01",X"EA",X"4E",X"64",X"00",X"D6",X"01",X"95",X"57",X"78",X"00",
		X"30",X"02",X"BF",X"59",X"46",X"00",X"62",X"02",X"BF",X"4C",X"28",X"00",X"00",X"FF",X"D8",X"09",
		X"00",X"00",X"03",X"FA",X"00",X"01",X"48",X"18",X"02",X"09",X"01",X"00",X"00",X"00",X"00",X"3F",
		X"90",X"01",X"00",X"00",X"00",X"3C",X"90",X"01",X"00",X"00",X"00",X"3D",X"90",X"01",X"18",X"00",
		X"00",X"3A",X"90",X"01",X"00",X"FF",X"30",X"09",X"DE",X"20",X"01",X"74",X"00",X"00",X"18",X"0A",
		X"04",X"0A",X"01",X"00",X"00",X"00",X"62",X"59",X"0A",X"00",X"1E",X"00",X"20",X"53",X"3C",X"00",
		X"1E",X"00",X"A1",X"55",X"1E",X"00",X"5A",X"00",X"E2",X"5B",X"28",X"00",X"64",X"00",X"62",X"59",
		X"1E",X"00",X"96",X"00",X"20",X"53",X"28",X"00",X"96",X"00",X"A1",X"55",X"32",X"00",X"BE",X"00",
		X"62",X"59",X"28",X"00",X"BE",X"00",X"E2",X"5B",X"28",X"00",X"00",X"FF",X"48",X"03",X"08",X"21",
		X"01",X"64",X"00",X"00",X"54",X"0A",X"01",X"01",X"04",X"0A",X"01",X"00",X"00",X"00",X"5F",X"4A",
		X"32",X"00",X"00",X"00",X"E0",X"51",X"32",X"00",X"0A",X"00",X"DF",X"4C",X"32",X"00",X"0A",X"00",
		X"60",X"4F",X"32",X"00",X"00",X"FF",X"D4",X"03",X"00",X"00",X"01",X"9E",X"00",X"00",X"04",X"0A",
		X"01",X"00",X"00",X"00",X"5F",X"4A",X"36",X"00",X"00",X"00",X"DF",X"4C",X"36",X"00",X"00",X"FF",
		X"EC",X"04",X"00",X"00",X"01",X"77",X"02",X"00",X"34",X"0A",X"05",X"14",X"01",X"0A",X"01",X"0B",
		X"00",X"00",X"08",X"0C",X"64",X"00",X"00",X"FF",X"1C",X"02",X"00",X"00",X"05",X"00",X"00",X"00",
		X"68",X"0A",X"02",X"DB",X"04",X"05",X"01",X"00",X"00",X"00",X"00",X"2E",X"2A",X"00",X"00",X"FF",
		X"80",X"02",X"00",X"00",X"06",X"60",X"01",X"00",X"58",X"0C",X"02",X"07",X"01",X"1E",X"02",X"51",
		X"00",X"00",X"00",X"2F",X"24",X"00",X"00",X"FF",X"78",X"03",X"00",X"00",X"02",X"39",X"01",X"00",
		X"08",X"0A",X"01",X"00",X"00",X"00",X"AA",X"31",X"0A",X"00",X"0A",X"00",X"B9",X"40",X"0A",X"00",
		X"14",X"00",X"05",X"4C",X"0A",X"00",X"00",X"FF",X"6B",X"03",X"00",X"00",X"14",X"70",X"00",X"FF",
		X"88",X"0D",X"04",X"00",X"01",X"00",X"00",X"00",X"00",X"36",X"28",X"00",X"0A",X"00",X"00",X"1E",
		X"32",X"00",X"B4",X"00",X"00",X"22",X"1E",X"00",X"B4",X"00",X"00",X"25",X"1E",X"00",X"B4",X"00",
		X"00",X"42",X"28",X"00",X"68",X"01",X"00",X"19",X"3C",X"00",X"EA",X"01",X"00",X"41",X"32",X"00",
		X"30",X"02",X"00",X"41",X"14",X"00",X"3A",X"02",X"00",X"25",X"3C",X"00",X"3A",X"02",X"00",X"3F",
		X"3C",X"00",X"44",X"02",X"00",X"22",X"28",X"00",X"A8",X"02",X"00",X"3D",X"3C",X"00",X"EE",X"02",
		X"00",X"3F",X"D2",X"00",X"F8",X"02",X"00",X"1E",X"6E",X"00",X"AC",X"03",X"00",X"22",X"32",X"00",
		X"AC",X"03",X"00",X"25",X"32",X"00",X"AC",X"03",X"00",X"3D",X"6E",X"00",X"10",X"04",X"00",X"3A",
		X"B4",X"00",X"6A",X"04",X"00",X"19",X"82",X"00",X"CE",X"04",X"00",X"3B",X"64",X"00",X"1E",X"05",
		X"00",X"22",X"32",X"00",X"1E",X"05",X"00",X"25",X"32",X"00",X"1E",X"05",X"00",X"3D",X"3C",X"00",
		X"E6",X"05",X"00",X"1D",X"28",X"00",X"E6",X"05",X"00",X"3F",X"A0",X"00",X"A4",X"06",X"00",X"3D",
		X"64",X"00",X"AE",X"06",X"00",X"20",X"32",X"00",X"AE",X"06",X"00",X"25",X"32",X"00",X"6C",X"07",
		X"00",X"19",X"A0",X"00",X"6C",X"07",X"00",X"3B",X"5A",X"00",X"D0",X"07",X"00",X"38",X"3C",X"00",
		X"34",X"08",X"00",X"20",X"3C",X"00",X"34",X"08",X"00",X"25",X"3C",X"00",X"A2",X"08",X"00",X"3D",
		X"32",X"00",X"F2",X"08",X"00",X"3F",X"B4",X"00",X"FC",X"08",X"00",X"1E",X"5A",X"00",X"B0",X"09",
		X"00",X"22",X"28",X"00",X"B0",X"09",X"00",X"25",X"28",X"00",X"BA",X"09",X"00",X"3D",X"3C",X"00",
		X"28",X"0A",X"00",X"3A",X"78",X"00",X"78",X"0A",X"00",X"19",X"A0",X"00",X"0E",X"0B",X"00",X"38",
		X"32",X"00",X"54",X"0B",X"00",X"22",X"46",X"00",X"5E",X"0B",X"00",X"25",X"32",X"00",X"68",X"0B",
		X"00",X"36",X"32",X"00",X"12",X"0C",X"00",X"1E",X"5A",X"00",X"12",X"0C",X"00",X"36",X"32",X"00",
		X"DA",X"0C",X"00",X"22",X"32",X"00",X"DA",X"0C",X"00",X"25",X"1E",X"00",X"DA",X"0C",X"00",X"42",
		X"6E",X"00",X"A2",X"0D",X"00",X"19",X"3C",X"00",X"10",X"0E",X"00",X"41",X"0A",X"00",X"60",X"0E",
		X"00",X"3F",X"64",X"00",X"6A",X"0E",X"00",X"22",X"3C",X"00",X"6A",X"0E",X"00",X"25",X"3C",X"00",
		X"6A",X"0E",X"00",X"41",X"14",X"00",X"CE",X"0E",X"00",X"3D",X"50",X"00",X"28",X"0F",X"00",X"1E",
		X"5A",X"00",X"28",X"0F",X"00",X"3F",X"D2",X"00",X"E6",X"0F",X"00",X"22",X"6E",X"00",X"E6",X"0F",
		X"00",X"25",X"46",X"00",X"F0",X"0F",X"00",X"3D",X"5A",X"00",X"54",X"10",X"00",X"3A",X"A0",X"00",
		X"86",X"10",X"00",X"19",X"AA",X"00",X"08",X"11",X"00",X"3B",X"64",X"00",X"58",X"11",X"00",X"22",
		X"3C",X"00",X"58",X"11",X"00",X"25",X"3C",X"00",X"58",X"11",X"00",X"3D",X"6E",X"00",X"20",X"12",
		X"00",X"3F",X"C8",X"00",X"2A",X"12",X"00",X"1D",X"46",X"00",X"E8",X"12",X"00",X"3D",X"BE",X"00",
		X"F2",X"12",X"00",X"20",X"46",X"00",X"F2",X"12",X"00",X"25",X"32",X"00",X"92",X"13",X"00",X"3B",
		X"78",X"00",X"B0",X"13",X"00",X"19",X"BE",X"00",X"1E",X"14",X"00",X"3A",X"32",X"00",X"64",X"14",
		X"00",X"38",X"32",X"00",X"6E",X"14",X"00",X"20",X"3C",X"00",X"78",X"14",X"00",X"25",X"3C",X"00",
		X"22",X"15",X"00",X"1E",X"64",X"00",X"2C",X"15",X"00",X"36",X"3C",X"00",X"EA",X"15",X"00",X"22",
		X"32",X"00",X"EA",X"15",X"00",X"25",X"1E",X"00",X"EA",X"15",X"00",X"3A",X"46",X"00",X"58",X"16",
		X"00",X"36",X"50",X"00",X"A8",X"16",X"00",X"19",X"BE",X"00",X"66",X"17",X"00",X"25",X"32",X"00",
		X"70",X"17",X"00",X"22",X"28",X"00",X"00",X"FF",X"48",X"18",X"DC",X"24",X"14",X"86",X"00",X"FF",
		X"C8",X"0B",X"09",X"0B",X"07",X"6E",X"01",X"00",X"00",X"00",X"00",X"0D",X"2D",X"00",X"BE",X"00",
		X"00",X"19",X"2D",X"00",X"18",X"01",X"00",X"0D",X"2D",X"00",X"7C",X"01",X"00",X"0D",X"2D",X"00",
		X"44",X"02",X"00",X"19",X"2D",X"00",X"A8",X"02",X"00",X"0D",X"2D",X"00",X"70",X"03",X"00",X"0D",
		X"2D",X"00",X"C0",X"03",X"00",X"19",X"2D",X"00",X"1A",X"04",X"00",X"0D",X"2D",X"00",X"7E",X"04",
		X"00",X"0D",X"2D",X"00",X"D8",X"04",X"00",X"0D",X"2D",X"00",X"46",X"05",X"00",X"19",X"2D",X"00",
		X"18",X"06",X"00",X"12",X"2D",X"00",X"CC",X"06",X"00",X"1E",X"2D",X"00",X"30",X"07",X"00",X"12",
		X"2D",X"00",X"94",X"07",X"00",X"12",X"2D",X"00",X"52",X"08",X"00",X"1E",X"2D",X"00",X"AC",X"08",
		X"00",X"12",X"2D",X"00",X"7E",X"09",X"00",X"12",X"2D",X"00",X"C4",X"09",X"00",X"1E",X"2D",X"00",
		X"28",X"0A",X"00",X"12",X"2D",X"00",X"8C",X"0A",X"00",X"12",X"2D",X"00",X"E6",X"0A",X"00",X"12",
		X"2D",X"00",X"40",X"0B",X"00",X"1E",X"2D",X"00",X"08",X"0C",X"00",X"14",X"2D",X"00",X"C6",X"0C",
		X"00",X"20",X"2D",X"00",X"20",X"0D",X"00",X"14",X"2D",X"00",X"8E",X"0D",X"00",X"14",X"2D",X"00",
		X"4C",X"0E",X"00",X"20",X"2D",X"00",X"B0",X"0E",X"00",X"14",X"2D",X"00",X"6E",X"0F",X"00",X"14",
		X"2D",X"00",X"C8",X"0F",X"00",X"20",X"2D",X"00",X"36",X"10",X"00",X"14",X"2D",X"00",X"90",X"10",
		X"00",X"14",X"2D",X"00",X"EA",X"10",X"00",X"14",X"2D",X"00",X"4E",X"11",X"00",X"20",X"2D",X"00",
		X"34",X"12",X"00",X"0D",X"2D",X"00",X"F2",X"12",X"00",X"19",X"2D",X"00",X"56",X"13",X"00",X"0D",
		X"2D",X"00",X"C4",X"13",X"00",X"0D",X"2D",X"00",X"78",X"14",X"00",X"19",X"2D",X"00",X"E6",X"14",
		X"00",X"0D",X"2D",X"00",X"9A",X"15",X"00",X"0D",X"2D",X"00",X"F4",X"15",X"00",X"19",X"2D",X"00",
		X"44",X"16",X"00",X"0D",X"2D",X"00",X"B2",X"16",X"00",X"0D",X"2D",X"00",X"20",X"17",X"00",X"0D",
		X"2D",X"00",X"70",X"17",X"00",X"19",X"2D",X"00",X"00",X"FF",X"3C",X"18",X"00",X"00",X"14",X"D4",
		X"00",X"FF",X"C8",X"0B",X"04",X"0B",X"07",X"6E",X"01",X"00",X"00",X"00",X"00",X"31",X"2D",X"00",
		X"B0",X"00",X"00",X"3D",X"2D",X"00",X"13",X"01",X"00",X"36",X"2D",X"00",X"81",X"01",X"00",X"38",
		X"2D",X"00",X"3C",X"02",X"00",X"3D",X"2D",X"00",X"9F",X"02",X"00",X"31",X"2D",X"00",X"5A",X"03",
		X"00",X"31",X"2D",X"00",X"BD",X"03",X"00",X"3D",X"2D",X"00",X"20",X"04",X"00",X"36",X"2D",X"00",
		X"83",X"04",X"00",X"38",X"2D",X"00",X"3E",X"05",X"00",X"3D",X"2D",X"00",X"F9",X"05",X"00",X"33",
		X"2D",X"00",X"BF",X"06",X"00",X"3F",X"2D",X"00",X"0C",X"07",X"00",X"38",X"2D",X"00",X"85",X"07",
		X"00",X"3A",X"2D",X"00",X"4B",X"08",X"00",X"3F",X"2D",X"00",X"B9",X"08",X"00",X"33",X"2D",X"00",
		X"74",X"09",X"00",X"33",X"2D",X"00",X"C1",X"09",X"00",X"3F",X"2D",X"00",X"24",X"0A",X"00",X"38",
		X"2D",X"00",X"92",X"0A",X"00",X"3A",X"2D",X"00",X"2C",X"0B",X"00",X"3F",X"2D",X"00",X"FD",X"0B",
		X"00",X"33",X"2D",X"00",X"B8",X"0C",X"00",X"36",X"2D",X"00",X"26",X"0D",X"00",X"38",X"2D",X"00",
		X"7E",X"0D",X"00",X"3D",X"2D",X"00",X"4F",X"0E",X"00",X"36",X"2D",X"00",X"B2",X"0E",X"00",X"38",
		X"2D",X"00",X"6D",X"0F",X"00",X"38",X"2D",X"00",X"DB",X"0F",X"00",X"3D",X"2D",X"00",X"96",X"10",
		X"00",X"36",X"2D",X"00",X"F9",X"10",X"00",X"38",X"2D",X"00",X"46",X"11",X"00",X"3D",X"2D",X"00",
		X"0C",X"12",X"00",X"31",X"2D",X"00",X"D2",X"12",X"00",X"36",X"2D",X"00",X"40",X"13",X"00",X"38",
		X"2D",X"00",X"98",X"13",X"00",X"3D",X"2D",X"00",X"5E",X"14",X"00",X"38",X"2D",X"00",X"E2",X"14",
		X"00",X"36",X"2D",X"00",X"92",X"15",X"00",X"3D",X"2D",X"00",X"00",X"16",X"00",X"38",X"2D",X"00",
		X"BB",X"16",X"00",X"36",X"2D",X"00",X"1E",X"17",X"00",X"31",X"2D",X"00",X"8C",X"17",X"00",X"36",
		X"2D",X"00",X"00",X"FF",X"3C",X"18",X"00",X"00",X"14",X"64",X"00",X"FF",X"C8",X"09",X"04",X"0B",
		X"07",X"C8",X"01",X"00",X"00",X"00",X"00",X"35",X"2D",X"00",X"05",X"00",X"00",X"19",X"2D",X"00",
		X"64",X"00",X"00",X"34",X"2D",X"00",X"91",X"00",X"00",X"20",X"2D",X"00",X"91",X"00",X"00",X"35",
		X"2D",X"00",X"F5",X"00",X"00",X"36",X"2D",X"00",X"27",X"01",X"00",X"22",X"2D",X"00",X"77",X"01",
		X"00",X"35",X"2D",X"00",X"AE",X"01",X"00",X"20",X"2D",X"00",X"AE",X"01",X"00",X"31",X"2D",X"00",
		X"0D",X"02",X"00",X"33",X"2D",X"00",X"35",X"02",X"00",X"19",X"2D",X"00",X"35",X"02",X"00",X"35",
		X"2D",X"00",X"94",X"02",X"00",X"34",X"2D",X"00",X"C6",X"02",X"00",X"35",X"2D",X"00",X"CB",X"02",
		X"00",X"20",X"2D",X"00",X"25",X"03",X"00",X"36",X"2D",X"00",X"4D",X"03",X"00",X"22",X"2D",X"00",
		X"A7",X"03",X"00",X"35",X"2D",X"00",X"D9",X"03",X"00",X"20",X"2D",X"00",X"D9",X"03",X"00",X"31",
		X"2D",X"00",X"38",X"04",X"00",X"33",X"2D",X"00",X"60",X"04",X"00",X"35",X"2D",X"00",X"65",X"04",
		X"00",X"19",X"2D",X"00",X"BF",X"04",X"00",X"34",X"2D",X"00",X"EC",X"04",X"00",X"20",X"2D",X"00",
		X"EC",X"04",X"00",X"35",X"2D",X"00",X"4B",X"05",X"00",X"36",X"2D",X"00",X"7D",X"05",X"00",X"22",
		X"2D",X"00",X"D7",X"05",X"00",X"35",X"2D",X"00",X"04",X"06",X"00",X"31",X"2D",X"00",X"09",X"06",
		X"00",X"20",X"2D",X"00",X"5E",X"06",X"00",X"33",X"2D",X"00",X"8B",X"06",X"00",X"35",X"2D",X"00",
		X"90",X"06",X"00",X"19",X"2D",X"00",X"0D",X"07",X"00",X"2C",X"2D",X"00",X"17",X"07",X"00",X"20",
		X"2D",X"00",X"6C",X"07",X"00",X"2E",X"2D",X"00",X"94",X"07",X"00",X"30",X"2D",X"00",X"A3",X"07",
		X"00",X"22",X"2D",X"00",X"EE",X"07",X"00",X"2E",X"2D",X"00",X"25",X"08",X"00",X"20",X"2D",X"00",
		X"2A",X"08",X"00",X"2C",X"2D",X"00",X"AC",X"08",X"00",X"14",X"2D",X"00",X"B1",X"08",X"00",X"33",
		X"2D",X"00",X"0B",X"09",X"00",X"32",X"2D",X"00",X"47",X"09",X"00",X"1B",X"2D",X"00",X"47",X"09",
		X"00",X"33",X"2D",X"00",X"9C",X"09",X"00",X"35",X"2D",X"00",X"C9",X"09",X"00",X"1D",X"2D",X"00",
		X"1E",X"0A",X"00",X"33",X"2D",X"00",X"50",X"0A",X"00",X"1B",X"2D",X"00",X"50",X"0A",X"00",X"30",
		X"2D",X"00",X"B4",X"0A",X"00",X"31",X"2D",X"00",X"D7",X"0A",X"00",X"14",X"2D",X"00",X"D7",X"0A",
		X"00",X"33",X"2D",X"00",X"36",X"0B",X"00",X"32",X"2D",X"00",X"63",X"0B",X"00",X"1B",X"2D",X"00",
		X"63",X"0B",X"00",X"33",X"2D",X"00",X"CC",X"0B",X"00",X"35",X"2D",X"00",X"FE",X"0B",X"00",X"1D",
		X"2D",X"00",X"49",X"0C",X"00",X"33",X"2D",X"00",X"7B",X"0C",X"00",X"30",X"2D",X"00",X"80",X"0C",
		X"00",X"1B",X"2D",X"00",X"D5",X"0C",X"00",X"31",X"2D",X"00",X"07",X"0D",X"00",X"33",X"2D",X"00",
		X"0C",X"0D",X"00",X"14",X"2D",X"00",X"6B",X"0D",X"00",X"32",X"2D",X"00",X"8E",X"0D",X"00",X"1B",
		X"2D",X"00",X"93",X"0D",X"00",X"33",X"2D",X"00",X"F2",X"0D",X"00",X"35",X"2D",X"00",X"2E",X"0E",
		X"00",X"1D",X"2D",X"00",X"7E",X"0E",X"00",X"33",X"2D",X"00",X"AB",X"0E",X"00",X"1B",X"2D",X"00",
		X"AB",X"0E",X"00",X"30",X"2D",X"00",X"05",X"0F",X"00",X"31",X"2D",X"00",X"37",X"0F",X"00",X"14",
		X"2D",X"00",X"37",X"0F",X"00",X"33",X"2D",X"00",X"BE",X"0F",X"00",X"2C",X"2D",X"00",X"C3",X"0F",
		X"00",X"1B",X"2D",X"00",X"18",X"10",X"00",X"2E",X"2D",X"00",X"45",X"10",X"00",X"30",X"2D",X"00",
		X"4A",X"10",X"00",X"1D",X"2D",X"00",X"9F",X"10",X"00",X"2E",X"2D",X"00",X"D1",X"10",X"00",X"1B",
		X"2D",X"00",X"D1",X"10",X"00",X"2C",X"2D",X"00",X"67",X"11",X"00",X"35",X"2D",X"00",X"6C",X"11",
		X"00",X"19",X"2D",X"00",X"C6",X"11",X"00",X"34",X"2D",X"00",X"F8",X"11",X"00",X"35",X"2D",X"00",
		X"FD",X"11",X"00",X"20",X"2D",X"00",X"57",X"12",X"00",X"36",X"2D",X"00",X"84",X"12",X"00",X"22",
		X"2D",X"00",X"DE",X"12",X"00",X"35",X"2D",X"00",X"0B",X"13",X"00",X"31",X"2D",X"00",X"10",X"13",
		X"00",X"20",X"2D",X"00",X"6A",X"13",X"00",X"33",X"2D",X"00",X"83",X"13",X"00",X"20",X"2D",X"00",
		X"97",X"13",X"00",X"35",X"2D",X"00",X"9C",X"13",X"00",X"19",X"2D",X"00",X"FB",X"13",X"00",X"34",
		X"2D",X"00",X"23",X"14",X"00",X"35",X"2D",X"00",X"28",X"14",X"00",X"20",X"2D",X"00",X"82",X"14",
		X"00",X"36",X"2D",X"00",X"B4",X"14",X"00",X"22",X"2D",X"00",X"04",X"15",X"00",X"35",X"2D",X"00",
		X"31",X"15",X"00",X"31",X"2D",X"00",X"36",X"15",X"00",X"20",X"2D",X"00",X"90",X"15",X"00",X"33",
		X"2D",X"00",X"C2",X"15",X"00",X"19",X"2D",X"00",X"C2",X"15",X"00",X"35",X"2D",X"00",X"21",X"16",
		X"00",X"34",X"2D",X"00",X"4E",X"16",X"00",X"35",X"2D",X"00",X"58",X"16",X"00",X"20",X"2D",X"00",
		X"AD",X"16",X"00",X"36",X"2D",X"00",X"E9",X"16",X"00",X"22",X"2D",X"00",X"39",X"17",X"00",X"35",
		X"2D",X"00",X"6B",X"17",X"00",X"20",X"2D",X"00",X"6B",X"17",X"00",X"31",X"2D",X"00",X"C0",X"17",
		X"00",X"33",X"2D",X"00",X"F2",X"17",X"00",X"35",X"2D",X"00",X"F7",X"17",X"00",X"19",X"2D",X"00",
		X"79",X"18",X"00",X"20",X"2D",X"00",X"79",X"18",X"00",X"2C",X"2D",X"00",X"D3",X"18",X"00",X"2E",
		X"2D",X"00",X"FB",X"18",X"00",X"30",X"2D",X"00",X"05",X"19",X"00",X"22",X"2D",X"00",X"5A",X"19",
		X"00",X"2E",X"2D",X"00",X"82",X"19",X"00",X"2C",X"2D",X"00",X"8C",X"19",X"00",X"20",X"2D",X"00",
		X"18",X"1A",X"00",X"1E",X"2D",X"00",X"18",X"1A",X"00",X"3A",X"2D",X"00",X"72",X"1A",X"00",X"39",
		X"2D",X"00",X"9F",X"1A",X"00",X"25",X"2D",X"00",X"9F",X"1A",X"00",X"3A",X"2D",X"00",X"F9",X"1A",
		X"00",X"3D",X"2D",X"00",X"30",X"1B",X"00",X"27",X"2D",X"00",X"7B",X"1B",X"00",X"3C",X"2D",X"00",
		X"AD",X"1B",X"00",X"3A",X"2D",X"00",X"B2",X"1B",X"00",X"25",X"2D",X"00",X"07",X"1C",X"00",X"38",
		X"2D",X"00",X"39",X"1C",X"00",X"1D",X"2D",X"00",X"39",X"1C",X"00",X"38",X"2D",X"00",X"A2",X"1C",
		X"00",X"37",X"2D",X"00",X"BB",X"1C",X"00",X"24",X"2D",X"00",X"CA",X"1C",X"00",X"38",X"2D",X"00",
		X"24",X"1D",X"00",X"3A",X"2D",X"00",X"56",X"1D",X"00",X"25",X"2D",X"00",X"A1",X"1D",X"00",X"38",
		X"2D",X"00",X"D3",X"1D",X"00",X"24",X"2D",X"00",X"D8",X"1D",X"00",X"36",X"2D",X"00",X"28",X"1E",
		X"00",X"35",X"2D",X"00",X"5F",X"1E",X"00",X"1B",X"2D",X"00",X"64",X"1E",X"00",X"35",X"2D",X"00",
		X"BE",X"1E",X"00",X"36",X"2D",X"00",X"EB",X"1E",X"00",X"22",X"2D",X"00",X"EB",X"1E",X"00",X"35",
		X"2D",X"00",X"40",X"1F",X"00",X"33",X"2D",X"00",X"86",X"1F",X"00",X"24",X"2D",X"00",X"D1",X"1F",
		X"00",X"31",X"2D",X"00",X"03",X"20",X"00",X"33",X"2D",X"00",X"08",X"20",X"00",X"22",X"2D",X"00",
		X"62",X"20",X"00",X"31",X"2D",X"00",X"94",X"20",X"00",X"19",X"2D",X"00",X"16",X"21",X"00",X"20",
		X"2D",X"00",X"9D",X"21",X"00",X"22",X"2D",X"00",X"29",X"22",X"00",X"20",X"2D",X"00",X"00",X"FF",
		X"B0",X"22",X"00",X"00",X"01",X"00",X"00",X"00",X"94",X"12",X"01",X"3B",X"02",X"0F",X"01",X"00",
		X"00",X"00",X"00",X"2C",X"99",X"00",X"00",X"FF",X"B2",X"02",X"00",X"00",X"01",X"00",X"00",X"00",
		X"94",X"0A",X"07",X"05",X"01",X"B8",X"01",X"00",X"00",X"00",X"00",X"2A",X"3C",X"00",X"00",X"FF",
		X"B2",X"02",X"38",X"2A",X"03",X"3A",X"02",X"00",X"14",X"0A",X"04",X"10",X"01",X"12",X"00",X"00",
		X"00",X"2C",X"14",X"00",X"00",X"FF",X"44",X"02",X"00",X"00",X"03",X"00",X"00",X"00",X"B4",X"0A",
		X"01",X"15",X"02",X"0A",X"02",X"10",X"02",X"12",X"28",X"00",X"00",X"29",X"96",X"00",X"00",X"FF",
		X"30",X"02",X"00",X"00",X"03",X"28",X"00",X"00",X"94",X"0A",X"02",X"01",X"04",X"2E",X"01",X"00",
		X"00",X"00",X"00",X"19",X"17",X"01",X"00",X"00",X"00",X"1E",X"17",X"01",X"00",X"00",X"00",X"20",
		X"17",X"01",X"0A",X"00",X"00",X"1B",X"17",X"01",X"0A",X"00",X"00",X"1D",X"17",X"01",X"0A",X"00",
		X"00",X"22",X"17",X"01",X"00",X"FF",X"FA",X"0A",X"00",X"00",X"01",X"5E",X"00",X"00",X"08",X"14",
		X"01",X"00",X"00",X"00",X"00",X"3D",X"55",X"00",X"05",X"00",X"00",X"22",X"46",X"00",X"0A",X"00",
		X"00",X"25",X"46",X"00",X"09",X"01",X"00",X"22",X"5A",X"00",X"09",X"01",X"00",X"3A",X"69",X"00",
		X"0E",X"01",X"00",X"1D",X"4B",X"00",X"0D",X"02",X"00",X"38",X"3C",X"00",X"0D",X"02",X"00",X"1D",
		X"2D",X"00",X"0D",X"02",X"00",X"20",X"28",X"00",X"25",X"03",X"00",X"1E",X"2D",X"00",X"2A",X"03",
		X"00",X"19",X"28",X"00",X"2A",X"03",X"00",X"36",X"28",X"00",X"2E",X"04",X"00",X"19",X"7D",X"00",
		X"2E",X"04",X"00",X"1D",X"82",X"00",X"33",X"04",X"00",X"35",X"7D",X"00",X"00",X"FF",X"7E",X"0E",
		X"46",X"2B",X"02",X"B6",X"00",X"00",X"08",X"0A",X"01",X"00",X"00",X"00",X"00",X"2E",X"64",X"00",
		X"14",X"00",X"00",X"1E",X"28",X"00",X"14",X"00",X"00",X"12",X"32",X"00",X"DC",X"00",X"00",X"11",
		X"3C",X"00",X"DC",X"00",X"00",X"2A",X"5A",X"00",X"E6",X"00",X"00",X"1D",X"28",X"00",X"4A",X"01",
		X"00",X"27",X"3C",X"00",X"54",X"01",X"00",X"0F",X"28",X"00",X"54",X"01",X"00",X"1B",X"28",X"00",
		X"44",X"02",X"00",X"0D",X"3C",X"00",X"44",X"02",X"00",X"19",X"3C",X"00",X"4E",X"02",X"00",X"25",
		X"5A",X"00",X"00",X"FF",X"78",X"0A",X"00",X"00",X"02",X"B6",X"00",X"00",X"08",X"0A",X"01",X"00",
		X"00",X"00",X"00",X"3A",X"68",X"01",X"DC",X"00",X"00",X"36",X"8C",X"00",X"54",X"01",X"00",X"33",
		X"18",X"01",X"4E",X"02",X"00",X"31",X"D2",X"00",X"00",X"FF",X"48",X"03",X"00",X"00",X"03",X"5E",
		X"00",X"00",X"08",X"1E",X"01",X"00",X"00",X"00",X"D5",X"59",X"42",X"00",X"8A",X"00",X"EF",X"57",
		X"30",X"00",X"0E",X"01",X"AA",X"56",X"36",X"00",X"98",X"01",X"C4",X"54",X"54",X"00",X"22",X"02",
		X"3C",X"52",X"54",X"00",X"A0",X"02",X"80",X"53",X"30",X"00",X"4E",X"03",X"C4",X"54",X"30",X"00",
		X"D2",X"03",X"66",X"55",X"42",X"00",X"5C",X"04",X"3C",X"52",X"30",X"00",X"00",X"FF",X"18",X"06",
		X"00",X"00",X"02",X"55",X"00",X"00",X"08",X"0E",X"01",X"00",X"00",X"00",X"00",X"3F",X"31",X"00",
		X"31",X"00",X"00",X"3D",X"23",X"00",X"62",X"00",X"00",X"3F",X"23",X"00",X"85",X"00",X"00",X"3D",
		X"2A",X"00",X"B6",X"00",X"00",X"3F",X"31",X"00",X"E0",X"00",X"00",X"3D",X"31",X"00",X"11",X"01",
		X"00",X"3F",X"38",X"00",X"42",X"01",X"00",X"3D",X"38",X"00",X"73",X"01",X"00",X"3F",X"38",X"00",
		X"A4",X"01",X"00",X"3D",X"5B",X"00",X"00",X"FF",X"17",X"03",X"00",X"00",X"02",X"00",X"00",X"FF",
		X"E8",X"13",X"07",X"24",X"04",X"0D",X"03",X"F8",X"01",X"05",X"00",X"00",X"00",X"31",X"10",X"01",
		X"00",X"FF",X"ED",X"03",X"C2",X"2D",X"03",X"6E",X"00",X"00",X"88",X"0C",X"09",X"00",X"01",X"00",
		X"00",X"00",X"07",X"35",X"49",X"00",X"78",X"00",X"07",X"36",X"49",X"00",X"E8",X"00",X"07",X"38",
		X"49",X"00",X"68",X"01",X"07",X"3A",X"49",X"00",X"E0",X"03",X"07",X"3A",X"49",X"00",X"60",X"04",
		X"07",X"3C",X"49",X"00",X"E0",X"04",X"07",X"3D",X"49",X"00",X"50",X"05",X"07",X"3F",X"49",X"00",
		X"D0",X"05",X"07",X"3D",X"49",X"00",X"50",X"06",X"07",X"3D",X"49",X"00",X"C0",X"06",X"07",X"3C",
		X"49",X"00",X"48",X"07",X"07",X"3C",X"49",X"00",X"B8",X"07",X"07",X"3A",X"49",X"00",X"40",X"08",
		X"07",X"3A",X"49",X"00",X"A8",X"08",X"07",X"38",X"49",X"00",X"38",X"09",X"07",X"38",X"49",X"00",
		X"88",X"0B",X"07",X"35",X"49",X"00",X"10",X"0C",X"07",X"36",X"49",X"00",X"90",X"0C",X"07",X"38",
		X"49",X"00",X"10",X"0D",X"07",X"3A",X"49",X"00",X"A0",X"0F",X"07",X"3A",X"49",X"00",X"10",X"10",
		X"07",X"3C",X"49",X"00",X"80",X"10",X"07",X"3D",X"49",X"00",X"F8",X"10",X"07",X"3F",X"49",X"00",
		X"88",X"11",X"07",X"3D",X"49",X"00",X"00",X"12",X"07",X"3D",X"49",X"00",X"78",X"12",X"07",X"3C",
		X"49",X"00",X"00",X"13",X"07",X"3C",X"49",X"00",X"70",X"13",X"07",X"3A",X"49",X"00",X"F8",X"13",
		X"07",X"3A",X"49",X"00",X"60",X"14",X"07",X"38",X"49",X"00",X"D8",X"14",X"07",X"38",X"49",X"00",
		X"C8",X"15",X"07",X"41",X"49",X"00",X"48",X"16",X"07",X"41",X"49",X"00",X"50",X"17",X"07",X"41",
		X"49",X"00",X"B8",X"17",X"07",X"42",X"49",X"00",X"28",X"18",X"07",X"41",X"49",X"00",X"A8",X"18",
		X"07",X"41",X"49",X"00",X"18",X"19",X"07",X"3F",X"49",X"00",X"98",X"19",X"07",X"3F",X"49",X"00",
		X"E8",X"1A",X"07",X"3F",X"49",X"00",X"60",X"1B",X"07",X"41",X"49",X"00",X"D8",X"1B",X"07",X"42",
		X"49",X"00",X"60",X"1C",X"07",X"42",X"49",X"00",X"D0",X"1C",X"07",X"41",X"49",X"00",X"58",X"1D",
		X"07",X"41",X"49",X"00",X"D0",X"1E",X"07",X"41",X"49",X"00",X"48",X"1F",X"07",X"42",X"49",X"00",
		X"B0",X"1F",X"07",X"41",X"49",X"00",X"20",X"20",X"07",X"44",X"49",X"00",X"90",X"20",X"07",X"42",
		X"49",X"00",X"10",X"21",X"07",X"42",X"49",X"00",X"78",X"22",X"07",X"3F",X"49",X"00",X"F0",X"22",
		X"07",X"41",X"49",X"00",X"60",X"23",X"07",X"42",X"49",X"00",X"D0",X"23",X"07",X"42",X"49",X"00",
		X"40",X"24",X"07",X"41",X"49",X"00",X"C0",X"24",X"07",X"41",X"49",X"00",X"20",X"26",X"07",X"41",
		X"49",X"00",X"90",X"26",X"07",X"42",X"49",X"00",X"00",X"27",X"07",X"44",X"49",X"00",X"68",X"27",
		X"07",X"46",X"49",X"00",X"70",X"27",X"07",X"46",X"49",X"00",X"58",X"29",X"07",X"46",X"49",X"00",
		X"D0",X"29",X"07",X"44",X"49",X"00",X"70",X"2B",X"07",X"46",X"49",X"00",X"E8",X"2B",X"07",X"42",
		X"49",X"00",X"28",X"2C",X"07",X"3F",X"49",X"00",X"E0",X"2C",X"07",X"3D",X"49",X"00",X"00",X"FF",
		X"D0",X"31",X"EA",X"30",X"04",X"6E",X"00",X"00",X"88",X"0C",X"09",X"00",X"01",X"00",X"77",X"00",
		X"00",X"19",X"49",X"00",X"77",X"00",X"00",X"23",X"49",X"00",X"77",X"00",X"00",X"25",X"49",X"00",
		X"5E",X"01",X"00",X"1E",X"49",X"00",X"E3",X"01",X"00",X"22",X"49",X"00",X"E3",X"01",X"00",X"25",
		X"49",X"00",X"6F",X"02",X"00",X"19",X"49",X"00",X"ED",X"02",X"00",X"22",X"49",X"00",X"ED",X"02",
		X"00",X"25",X"49",X"00",X"79",X"03",X"00",X"1E",X"49",X"00",X"F0",X"03",X"00",X"25",X"49",X"00",
		X"F7",X"03",X"00",X"22",X"49",X"00",X"67",X"04",X"00",X"19",X"49",X"00",X"DE",X"04",X"00",X"22",
		X"49",X"00",X"E5",X"04",X"00",X"25",X"49",X"00",X"63",X"05",X"00",X"1E",X"49",X"00",X"DA",X"05",
		X"00",X"24",X"49",X"00",X"DA",X"05",X"00",X"27",X"49",X"00",X"58",X"06",X"00",X"1B",X"49",X"00",
		X"C8",X"06",X"00",X"24",X"49",X"00",X"C8",X"06",X"00",X"27",X"49",X"00",X"46",X"07",X"00",X"20",
		X"49",X"00",X"C4",X"07",X"00",X"24",X"49",X"00",X"C4",X"07",X"00",X"27",X"49",X"00",X"34",X"08",
		X"00",X"1B",X"49",X"00",X"B2",X"08",X"00",X"27",X"49",X"00",X"B9",X"08",X"00",X"24",X"49",X"00",
		X"29",X"09",X"00",X"1D",X"49",X"00",X"A0",X"09",X"00",X"20",X"49",X"00",X"A0",X"09",X"00",X"25",
		X"49",X"00",X"25",X"0A",X"00",X"19",X"49",X"00",X"9C",X"0A",X"00",X"20",X"49",X"00",X"9C",X"0A",
		X"00",X"25",X"49",X"00",X"1A",X"0B",X"00",X"1D",X"49",X"00",X"08",X"0C",X"00",X"19",X"49",X"00",
		X"08",X"0C",X"00",X"23",X"49",X"00",X"08",X"0C",X"00",X"25",X"49",X"00",X"12",X"0D",X"00",X"1E",
		X"49",X"00",X"89",X"0D",X"00",X"22",X"49",X"00",X"89",X"0D",X"00",X"25",X"49",X"00",X"0E",X"0E",
		X"00",X"19",X"49",X"00",X"8C",X"0E",X"00",X"22",X"49",X"00",X"8C",X"0E",X"00",X"25",X"49",X"00",
		X"11",X"0F",X"00",X"1E",X"49",X"00",X"88",X"0F",X"00",X"22",X"49",X"00",X"88",X"0F",X"00",X"25",
		X"49",X"00",X"1B",X"10",X"00",X"19",X"49",X"00",X"92",X"10",X"00",X"22",X"49",X"00",X"92",X"10",
		X"00",X"25",X"49",X"00",X"17",X"11",X"00",X"1E",X"49",X"00",X"79",X"11",X"00",X"24",X"49",X"00",
		X"80",X"11",X"00",X"27",X"49",X"00",X"05",X"12",X"00",X"1B",X"49",X"00",X"75",X"12",X"00",X"24",
		X"49",X"00",X"75",X"12",X"00",X"27",X"49",X"00",X"FA",X"12",X"00",X"20",X"49",X"00",X"6A",X"13",
		X"00",X"24",X"49",X"00",X"6A",X"13",X"00",X"27",X"49",X"00",X"EF",X"13",X"00",X"1B",X"49",X"00",
		X"58",X"14",X"00",X"27",X"49",X"00",X"66",X"14",X"00",X"24",X"49",X"00",X"DD",X"14",X"00",X"1D",
		X"49",X"00",X"54",X"15",X"00",X"20",X"49",X"00",X"5B",X"15",X"00",X"25",X"49",X"00",X"D9",X"15",
		X"00",X"19",X"49",X"00",X"49",X"16",X"00",X"25",X"49",X"00",X"50",X"16",X"00",X"20",X"49",X"00",
		X"C7",X"16",X"00",X"1D",X"49",X"00",X"45",X"17",X"00",X"20",X"49",X"00",X"45",X"17",X"00",X"25",
		X"49",X"00",X"C3",X"17",X"00",X"19",X"49",X"00",X"33",X"18",X"00",X"20",X"49",X"00",X"33",X"18",
		X"00",X"25",X"49",X"00",X"AA",X"18",X"00",X"1E",X"49",X"00",X"2F",X"19",X"00",X"23",X"49",X"00",
		X"2F",X"19",X"00",X"27",X"49",X"00",X"A6",X"19",X"00",X"1B",X"49",X"00",X"16",X"1A",X"00",X"23",
		X"49",X"00",X"1D",X"1A",X"00",X"27",X"49",X"00",X"55",X"1A",X"00",X"23",X"49",X"00",X"94",X"1A",
		X"00",X"1E",X"49",X"00",X"0B",X"1B",X"00",X"23",X"49",X"00",X"0B",X"1B",X"00",X"27",X"49",X"00",
		X"7B",X"1B",X"00",X"1B",X"49",X"00",X"E4",X"1B",X"00",X"23",X"49",X"00",X"F2",X"1B",X"00",X"27",
		X"49",X"00",X"70",X"1C",X"00",X"20",X"49",X"00",X"D9",X"1C",X"00",X"25",X"49",X"00",X"E0",X"1C",
		X"00",X"29",X"49",X"00",X"49",X"1D",X"00",X"1D",X"49",X"00",X"C7",X"1D",X"00",X"25",X"49",X"00",
		X"C7",X"1D",X"00",X"29",X"49",X"00",X"3E",X"1E",X"00",X"20",X"49",X"00",X"C3",X"1E",X"00",X"25",
		X"49",X"00",X"C3",X"1E",X"00",X"29",X"49",X"00",X"41",X"1F",X"00",X"1D",X"49",X"00",X"B8",X"1F",
		X"00",X"25",X"49",X"00",X"BF",X"1F",X"00",X"29",X"49",X"00",X"28",X"20",X"00",X"1E",X"49",X"00",
		X"9F",X"20",X"00",X"23",X"49",X"00",X"9F",X"20",X"00",X"27",X"49",X"00",X"16",X"21",X"00",X"1B",
		X"49",X"00",X"8D",X"21",X"00",X"23",X"49",X"00",X"94",X"21",X"00",X"27",X"49",X"00",X"04",X"22",
		X"00",X"1E",X"49",X"00",X"74",X"22",X"00",X"23",X"49",X"00",X"7B",X"22",X"00",X"27",X"49",X"00",
		X"EB",X"22",X"00",X"1B",X"49",X"00",X"5B",X"23",X"00",X"23",X"49",X"00",X"5B",X"23",X"00",X"27",
		X"49",X"00",X"D2",X"23",X"00",X"20",X"49",X"00",X"49",X"24",X"00",X"25",X"49",X"00",X"57",X"24",
		X"00",X"29",X"49",X"00",X"B9",X"24",X"00",X"1D",X"49",X"00",X"30",X"25",X"00",X"25",X"49",X"00",
		X"37",X"25",X"00",X"29",X"49",X"00",X"A0",X"25",X"00",X"20",X"49",X"00",X"17",X"26",X"00",X"25",
		X"49",X"00",X"1E",X"26",X"00",X"29",X"49",X"00",X"95",X"26",X"00",X"1D",X"49",X"00",X"FE",X"26",
		X"00",X"25",X"49",X"00",X"FE",X"26",X"00",X"29",X"49",X"00",X"91",X"27",X"00",X"1E",X"49",X"00",
		X"91",X"27",X"00",X"22",X"49",X"00",X"98",X"27",X"00",X"25",X"49",X"00",X"4A",X"29",X"00",X"20",
		X"49",X"00",X"4A",X"29",X"00",X"24",X"49",X"00",X"4A",X"29",X"00",X"27",X"49",X"00",X"3B",X"2B",
		X"00",X"22",X"49",X"00",X"D5",X"2B",X"00",X"1E",X"49",X"00",X"0D",X"2C",X"00",X"1B",X"49",X"00",
		X"D8",X"2C",X"00",X"19",X"49",X"00",X"00",X"FF",X"80",X"2D",X"00",X"00",X"04",X"6E",X"00",X"00",
		X"88",X"0C",X"09",X"00",X"01",X"00",X"81",X"01",X"00",X"12",X"49",X"00",X"6F",X"02",X"00",X"0D",
		X"49",X"00",X"79",X"03",X"00",X"12",X"49",X"00",X"67",X"04",X"00",X"0D",X"49",X"00",X"63",X"05",
		X"00",X"12",X"49",X"00",X"3C",X"06",X"00",X"0F",X"49",X"00",X"38",X"07",X"00",X"14",X"49",X"00",
		X"3B",X"08",X"00",X"0F",X"49",X"00",X"22",X"09",X"00",X"11",X"49",X"00",X"25",X"0A",X"00",X"0D",
		X"49",X"00",X"1A",X"0B",X"00",X"11",X"49",X"00",X"20",X"0D",X"00",X"12",X"49",X"00",X"23",X"0E",
		X"00",X"0D",X"49",X"00",X"1F",X"0F",X"00",X"12",X"49",X"00",X"1B",X"10",X"00",X"0D",X"49",X"00",
		X"09",X"11",X"00",X"12",X"49",X"00",X"FE",X"11",X"00",X"0F",X"49",X"00",X"08",X"13",X"00",X"14",
		X"49",X"00",X"FD",X"13",X"00",X"0F",X"49",X"00",X"EB",X"14",X"00",X"11",X"49",X"00",X"EE",X"15",
		X"00",X"0D",X"49",X"00",X"E3",X"16",X"00",X"11",X"49",X"00",X"BC",X"17",X"00",X"0D",X"49",X"00",
		X"B1",X"18",X"00",X"12",X"49",X"00",X"A6",X"19",X"00",X"0F",X"49",X"00",X"9B",X"1A",X"00",X"12",
		X"49",X"00",X"74",X"1B",X"00",X"0F",X"49",X"00",X"5B",X"1C",X"00",X"11",X"49",X"00",X"5E",X"1D",
		X"00",X"0D",X"49",X"00",X"61",X"1E",X"00",X"11",X"49",X"00",X"4F",X"1F",X"00",X"0D",X"49",X"00",
		X"2F",X"20",X"00",X"12",X"49",X"00",X"1D",X"21",X"00",X"0F",X"49",X"00",X"0B",X"22",X"00",X"12",
		X"49",X"00",X"F2",X"22",X"00",X"0F",X"49",X"00",X"D9",X"23",X"00",X"11",X"49",X"00",X"B9",X"24",
		X"00",X"0D",X"49",X"00",X"B5",X"25",X"00",X"11",X"49",X"00",X"9C",X"26",X"00",X"0D",X"49",X"00",
		X"8A",X"27",X"00",X"12",X"49",X"00",X"7B",X"29",X"00",X"14",X"49",X"00",X"00",X"FF",X"59",X"2E",
		X"00",X"00",X"03",X"CF",X"00",X"00",X"08",X"32",X"01",X"00",X"00",X"00",X"00",X"3D",X"36",X"00",
		X"06",X"00",X"00",X"36",X"30",X"00",X"06",X"00",X"00",X"38",X"30",X"00",X"EA",X"00",X"00",X"31",
		X"3C",X"00",X"F0",X"00",X"00",X"33",X"30",X"00",X"F0",X"00",X"00",X"38",X"36",X"00",X"E0",X"01",
		X"00",X"2E",X"42",X"00",X"E0",X"01",X"00",X"30",X"3C",X"00",X"E0",X"01",X"00",X"35",X"3C",X"00",
		X"EC",X"01",X"00",X"31",X"06",X"00",X"C4",X"02",X"00",X"2A",X"2A",X"00",X"C4",X"02",X"00",X"2C",
		X"2A",X"00",X"C4",X"02",X"00",X"31",X"2A",X"00",X"CC",X"03",X"00",X"2E",X"54",X"00",X"CC",X"03",
		X"00",X"30",X"54",X"00",X"CC",X"03",X"00",X"35",X"5A",X"00",X"00",X"FF",X"4E",X"06",X"00",X"00",
		X"02",X"7D",X"01",X"00",X"88",X"0A",X"01",X"D2",X"01",X"00",X"00",X"00",X"1C",X"4C",X"32",X"00",
		X"0A",X"00",X"97",X"4C",X"32",X"00",X"00",X"FF",X"D0",X"02",X"00",X"00",X"04",X"5F",X"00",X"00",
		X"C8",X"0A",X"0A",X"1A",X"06",X"FF",X"01",X"00",X"00",X"00",X"00",X"16",X"0F",X"04",X"1E",X"00",
		X"00",X"20",X"0F",X"04",X"1E",X"00",X"00",X"27",X"0F",X"04",X"28",X"00",X"00",X"29",X"0F",X"04",
		X"32",X"00",X"00",X"19",X"0F",X"04",X"3C",X"00",X"00",X"1B",X"0F",X"04",X"00",X"FF",X"08",X"07",
		X"00",X"00",X"03",X"02",X"02",X"00",X"48",X"0A",X"02",X"F0",X"01",X"00",X"00",X"00",X"F9",X"1B",
		X"69",X"00",X"00",X"FF",X"DA",X"02",X"00",X"00",X"03",X"90",X"01",X"00",X"68",X"0A",X"04",X"FA",
		X"02",X"0E",X"01",X"05",X"00",X"00",X"D9",X"0A",X"28",X"00",X"00",X"00",X"26",X"33",X"28",X"00",
		X"00",X"00",X"FF",X"3D",X"32",X"00",X"00",X"FF",X"A0",X"05",X"00",X"00",X"04",X"D6",X"01",X"00",
		X"68",X"0A",X"04",X"FA",X"02",X"0E",X"01",X"00",X"00",X"00",X"99",X"12",X"28",X"00",X"00",X"00",
		X"73",X"1D",X"28",X"00",X"00",X"FF",X"A8",X"02",X"00",X"00",X"03",X"00",X"00",X"00",X"E8",X"06",
		X"05",X"03",X"02",X"01",X"03",X"30",X"01",X"42",X"00",X"00",X"00",X"20",X"90",X"01",X"00",X"00",
		X"00",X"22",X"90",X"01",X"00",X"00",X"00",X"2E",X"90",X"01",X"00",X"FF",X"36",X"03",X"00",X"00",
		X"03",X"00",X"00",X"00",X"E8",X"06",X"05",X"03",X"05",X"01",X"03",X"30",X"01",X"42",X"00",X"00",
		X"BA",X"29",X"90",X"01",X"00",X"00",X"44",X"40",X"90",X"01",X"00",X"FF",X"08",X"04",X"80",X"33",
		X"03",X"00",X"00",X"00",X"E8",X"08",X"05",X"15",X"02",X"D5",X"03",X"5F",X"01",X"42",X"00",X"00",
		X"00",X"19",X"19",X"00",X"00",X"00",X"00",X"1C",X"19",X"00",X"12",X"00",X"00",X"20",X"19",X"00",
		X"12",X"00",X"00",X"27",X"19",X"00",X"1E",X"00",X"00",X"29",X"19",X"00",X"00",X"FF",X"78",X"03",
		X"00",X"00",X"03",X"B6",X"00",X"00",X"C8",X"0A",X"01",X"25",X"02",X"2A",X"01",X"00",X"6B",X"00",
		X"CF",X"4A",X"69",X"00",X"C5",X"00",X"F5",X"55",X"69",X"00",X"01",X"01",X"28",X"4D",X"69",X"00",
		X"6F",X"01",X"21",X"57",X"69",X"00",X"E7",X"01",X"F5",X"55",X"69",X"00",X"23",X"02",X"28",X"4D",
		X"69",X"00",X"AF",X"02",X"21",X"57",X"69",X"00",X"31",X"03",X"F5",X"55",X"69",X"00",X"00",X"FF",
		X"B4",X"0A",X"00",X"00",X"03",X"00",X"00",X"00",X"68",X"0A",X"06",X"20",X"03",X"73",X"01",X"03",
		X"00",X"00",X"00",X"2F",X"15",X"00",X"00",X"FF",X"31",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"68",X"0A",X"06",X"20",X"03",X"73",X"01",X"03",X"00",X"00",X"00",X"33",X"15",X"00",X"00",X"FF",
		X"4B",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"68",X"0A",X"06",X"20",X"03",X"73",X"01",X"03",
		X"00",X"00",X"00",X"3B",X"15",X"00",X"00",X"FF",X"6A",X"00",X"34",X"34",X"02",X"5F",X"01",X"00",
		X"C8",X"0A",X"09",X"01",X"09",X"F7",X"01",X"00",X"61",X"00",X"B3",X"15",X"7D",X"00",X"61",X"00",
		X"A6",X"23",X"7D",X"00",X"6B",X"00",X"26",X"33",X"7D",X"00",X"7F",X"00",X"BF",X"45",X"7D",X"00",
		X"00",X"FF",X"F4",X"06",X"00",X"00",X"02",X"74",X"00",X"00",X"14",X"08",X"04",X"0A",X"01",X"00",
		X"00",X"00",X"00",X"27",X"3C",X"00",X"1E",X"00",X"00",X"33",X"32",X"00",X"00",X"FF",X"0C",X"03",
		X"00",X"00",X"03",X"00",X"00",X"00",X"C8",X"06",X"09",X"FF",X"02",X"FD",X"02",X"47",X"00",X"00",
		X"00",X"20",X"31",X"00",X"00",X"FF",X"4A",X"01",X"00",X"00",X"03",X"00",X"00",X"00",X"C8",X"06",
		X"09",X"FF",X"02",X"FD",X"02",X"47",X"00",X"00",X"00",X"25",X"31",X"00",X"00",X"FF",X"A4",X"01",
		X"00",X"00",X"03",X"00",X"00",X"00",X"C8",X"06",X"09",X"FF",X"02",X"FD",X"02",X"47",X"00",X"00",
		X"00",X"2C",X"31",X"00",X"00",X"FF",X"F6",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"C8",X"06",
		X"09",X"FF",X"02",X"FD",X"02",X"47",X"00",X"00",X"00",X"30",X"31",X"00",X"00",X"FF",X"6E",X"01",
		X"00",X"00",X"03",X"00",X"00",X"00",X"C8",X"06",X"09",X"FF",X"02",X"FD",X"02",X"47",X"00",X"00",
		X"00",X"33",X"31",X"00",X"00",X"FF",X"10",X"02",X"00",X"00",X"03",X"00",X"00",X"00",X"C8",X"06",
		X"09",X"FF",X"02",X"FD",X"02",X"47",X"00",X"00",X"00",X"36",X"31",X"00",X"00",X"FF",X"F6",X"00",
		X"00",X"10",X"00",X"10",X"0E",X"10",X"40",X"10",X"DC",X"11",X"02",X"12",X"22",X"12",X"FE",X"17",
		X"60",X"1D",X"7A",X"1D",X"94",X"1D",X"AA",X"1D",X"C0",X"1D",X"D8",X"1D",X"F2",X"1D",X"3C",X"1E",
		X"5C",X"1E",X"72",X"1E",X"9E",X"1E",X"B6",X"1E",X"0A",X"1F",X"70",X"20",X"98",X"20",X"22",X"21",
		X"3A",X"21",X"52",X"21",X"00",X"10",X"00",X"10",X"6A",X"21",X"8A",X"21",X"AA",X"23",X"F6",X"25",
		X"F2",X"29",X"0A",X"2A",X"22",X"2A",X"52",X"2A",X"88",X"2A",X"F0",X"2A",X"6C",X"2B",X"B0",X"2B",
		X"FA",X"2B",X"14",X"2C",X"F0",X"31",X"5E",X"32",X"7A",X"32",X"B0",X"32",X"C6",X"32",X"EA",X"32",
		X"08",X"33",X"2E",X"33",X"4E",X"33",X"C2",X"33",X"DA",X"33",X"F2",X"33",X"0A",X"34",X"50",X"34",
		X"68",X"34",X"80",X"34",X"98",X"34",X"B0",X"34",X"C8",X"34",X"00",X"00",X"05",X"01",X"0C",X"02",
		X"19",X"03",X"27",X"04",X"32",X"05",X"62",X"08",X"8D",X"0B",X"D2",X"0F",X"FF",X"01",X"00",X"00",
		X"0A",X"0F",X"FF",X"0F",X"00",X"0A",X"FF",X"0A",X"00",X"0A",X"64",X"0F",X"A0",X"0F",X"FF",X"00",
		X"00",X"00",X"05",X"05",X"0F",X"0A",X"14",X"0C",X"19",X"0F",X"1B",X"0F",X"1E",X"0C",X"23",X"0A",
		X"28",X"05",X"41",X"03",X"64",X"01",X"FF",X"00",X"00",X"03",X"27",X"04",X"32",X"05",X"62",X"08",
		X"8D",X"0B",X"D2",X"0F",X"FF",X"00",X"00",X"0D",X"FF",X"0D",X"00",X"00",X"28",X"02",X"32",X"03",
		X"4B",X"07",X"5F",X"0D",X"6B",X"0E",X"73",X"0F",X"80",X"0E",X"9A",X"08",X"B8",X"04",X"FF",X"00",
		X"5A",X"35",X"6E",X"35",X"00",X"10",X"74",X"35",X"78",X"35",X"00",X"10",X"80",X"35",X"98",X"35",
		X"A6",X"35",X"AA",X"35",X"00",X"00",X"18",X"E0",X"FF",X"92",X"00",X"06",X"F1",X"FF",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"08",X"00",X"E2",X"70",X"07",X"92",X"00",X"FF",X"00",X"18",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"13",X"00",X"19",X"33",X"01",X"24",X"00",X"4B",X"66",X"08",
		X"43",X"00",X"7D",X"99",X"15",X"2B",X"00",X"84",X"CC",X"16",X"14",X"00",X"8D",X"85",X"17",X"0D",
		X"00",X"96",X"00",X"18",X"00",X"00",X"FF",X"00",X"18",X"00",X"00",X"00",X"3D",X"00",X"5A",X"99",
		X"15",X"3D",X"00",X"64",X"00",X"18",X"00",X"00",X"69",X"00",X"18",X"C2",X"FF",X"73",X"99",X"15",
		X"C2",X"FF",X"CD",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"16",X"00",X"FF",
		X"94",X"16",X"00",X"00",X"00",X"00",X"00",X"69",X"37",X"00",X"01",X"00",X"C8",X"DC",X"00",X"DF",
		X"FF",X"D2",X"92",X"FF",X"00",X"00",X"FF",X"92",X"FF",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"E7",X"FF",X"5A",X"0B",X"FF",X"DF",X"FF",X"5F",X"68",X"FE",X"3D",X"00",X"61",X"E2",X"FE",
		X"77",X"00",X"71",X"5D",X"06",X"03",X"00",X"A6",X"29",X"07",X"03",X"00",X"C1",X"8F",X"07",X"B7",
		X"FF",X"C8",X"91",X"05",X"4C",X"00",X"D0",X"F5",X"07",X"9A",X"FF",X"D6",X"91",X"05",X"55",X"00",
		X"DC",X"8F",X"07",X"D0",X"FF",X"EC",X"9D",X"04",X"76",X"00",X"F2",X"66",X"07",X"CD",X"FF",X"FA",
		X"CF",X"05",X"6E",X"00",X"FF",X"F5",X"07",X"D4",X"35",X"D4",X"35",X"E1",X"35",X"EE",X"35",X"19",
		X"36",X"3A",X"36",X"42",X"36",X"00",X"10",X"59",X"36",X"00",X"0F",X"05",X"08",X"64",X"00",X"9C",
		X"00",X"FA",X"08",X"FF",X"0F",X"00",X"0A",X"64",X"00",X"FF",X"06",X"00",X"03",X"00",X"03",X"FF",
		X"03",X"00",X"05",X"FF",X"0C",X"00",X"10",X"B9",X"36",X"C5",X"36",X"CB",X"36",X"D1",X"36",X"00",
		X"1E",X"FF",X"00",X"00",X"1F",X"FF",X"00",X"00",X"06",X"06",X"06",X"FF",X"06",X"00",X"09",X"00",
		X"09",X"FF",X"09",X"DF",X"36",X"E3",X"36",X"E7",X"36",X"ED",X"36",X"00",X"01",X"80",X"00",X"FF",
		X"00",X"FB",X"36",X"00",X"01",X"80",X"00",X"FF",X"00",X"03",X"37",X"00",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
